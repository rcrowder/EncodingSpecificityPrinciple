BZh91AY&SY�z���߀rp����� ����bh? |� "      H�n���@                                     />�E
Q%*���R�� ��!ET(��%TE*UER�UQP$B�U!缀	P%D�ETPPEJHIER���@���J�QB��T�$�U*�E 
*�PU�@l�y"A��R���p}� �ީ*��z�Xu 9�UgaЉ���A^�P��X;.^�2Wy���-��@���I�\t7XT=��URT�R�  
�HU�ʟ|�
>��{�� z�o>U��ϏE}�<|L ���OUm��P�ް{�.�7��{8<X��n�a&z�yJ���zR�DC�� TUIR����@S�H��w�"���D1O{�dw�Iz�&{��UW�=*����Мcu�9:p�Z��T���u"C�*����w�*sv�)ABT@�J�4��{�v�T�nyR;�;�*��c�3Zi��F6[j��7�R���D��J�s������2�8��3����*@TE�TPAJ�)T*)� ��T9�^ꔧ���ܫH��r���n���@c�QUo8󞲌���Ltk݃�����7�)TN�$����R��{<0j��tO%H$��QUB��I)'Vi1�Y�=�"�w��R��OTƚ{�:���7
O)g�q�U^]�Ep���{uzI�����F��R��c�c�Rz�U"�EࠩR�R�@��JR��)8g<���Cє{�OR1^���bg#J*�A�s�Jw3��a[�wDW�����To{uAQ�R,3���,�c��%��U*)H�*��޻�C�c��)A��<c�+�.��dVh�z��S{t�&rЩN�=*��wz
�8z��wA���<'��/Z2DUQD��JP(*�Q��P�8R�Y�����u�Hi�h8���C�r�N�@�f�������<A�`I���T�Uy�X���U��p�
P�H�"�R���^�������{ґq���� w6N7=�U'�Ǡ���Rq��*���י�95y�ް�                               SѠҔ�H�h�h A�  "��%*�� 40 i�0L=�$h��       i�T����	�� &  4уOHI�T�C i�M144i��d0L#@�����4L'�z�5=&�~���<&ҟO��'�W����w��u���y���o]z�n�=��2�����ΔUW�� �J*��J��E��"UW"���R��]�˟����?.������������EUgǍ��U���Z�Y��ve�ڝڪ����������._S���_�QC���u�v���~�����ݷ��ߛxg}�v�l�n������s�9˾m�.��v�3�l�;�g�+
��1}O�`�RF	X���XF�1I�TP�d�$X/͗�w�;g�u�]cf�X���=i���\\i��ƽk�<<kn�}x�g��c�������<���燝6:Ӷ��;��l۶<�9λk��z���x����3֝�ֽ�����k��8�δ��w�������sc������X.qŊ�v�ȡe6C$�
�a
�e�$^"E�(�H��.����s���_?]��B�����3�	11GE�(R`�D0����%$/��R|IH^���PĐ@(\<p�SR/
0A�&|)8+"�-x� 	����E`.��&Y�F
�B����b|�%�,���BI�X�/����<+돏Zyβ��v�wZ�=ns�[E�;k�y�<g�z�9ǝS�v�ym�.4^q�W�q��v�l��kƮt��DxP�%�(����Ł6�����D�Z�_J(���t����>���8�p	 (��4�$K��ڛ|
(\$��$��u�����Ӣg	(\(�ǅқ�ӂ��v���8�I�J��^�R��:��ָԽ��T���y�u�x�{�Wl�'9N��b�Ry�Ƃ�Q�s���ҹ��*�Ke]�/Y���q��Ҟ4G|/.2#���&���6�֋�N�z�s���b�2v��U�^�6Ch����*��	��iz�wձW|�jy��I�T:�:�zĽ�ʯ��I�)�S�S�T�*�<h:�zѴ��u��;�GY*���!�J4/�=꧝)�%ơzʹ�w�zʼ�{��C��XmK֫j���R��֗9YW��8���%Έ�;���=����+�/y.r��y��E���j6���zÍj��=i<���A�Ds��u��uS��u�s��(���ꇼ���hv��Jy�l��\iC�O9<�9�q��	�;�<d�:�yO:<�1l��Ʈu]�t���i6WYyҸ�s����]�/ZOxu�ު�:]�9��//Y�9���.�Oz�|N4<�x˶�z�.4��lr8�9��)��K���S�T�N��ꮵS�^��+�K���mT��S��q�����s��h�i=�z���9�iO��E�Sj�e;eNrN4�x���^�ļ`��֭�֥�����Nps��OY��Z^2N5�Jv�X�X/�2��zԽ�ʜ�e;h{��Q���dڻeU�#���T���Q�Q�%�I�^�������9�{�s�;eN�S���*v�{�6�mS�K�S���U�/z���l��l��OY^�z��u�{�u�X��Z��F�z��N�u�mrw���W�c��퇍)�Ce<�ڽ�=�2�`��u�m�G|�s�z��I֫�P�IG��8����v+0b����τ�,#������xBA:z�l�^��w��;e�/;�.��x��w�ۍw����z��vӍ��<��;c�ll{��:�|`�D��<Ց�I� @�.�t�:/��2��X,���"�#��a)G�gCV*0O�xRB ����X��	>�T.���R+,@�Q�	� ,,L��2 �;�<;�:������0�<�nsk���'�zͺ��w���o�/���N<o��$I6�?h?�W��&SRa�W�[P��I:��F�;����ѷ)��,�G3�F��*P]�T�a�.u�g��_r�n�د@G����=���q#�uKʡ�=��\ԓ���]��F�����E�_��6c`3�s���rs^E1�͹sĪ��p�fT=�վ�.��L��|���|��+��듕������ܚ�Vs^�H"Q����{�l�4�4y�;&���S����S��� ~V��2�Η��p����Nz�X���:E� �����+x�ou!m@k�n�[Wk�<��=���W*3�FE�=�X�>���
��d˫�0��f�U����+�&L�wk����r�����T���n���F�^��X|�8-<u��;��v^�S��Z �U��:ϻ���,rfۘ�ܢa{9h��B��,KG��t�ڣGՍ��%�s(�"��^nƽ���m϶�����ֽ�r�}�H��g�g�|�NJ��Y��<����;�0�&�]s�{5f}�
gg�+Z���I,�f�{j���n�P��M]�����-xX�Ќ(㰽��t��&���oX��i��=w-툘7q ^\����q�zI��w�HV�㼻��y����ɼ�l��C7����
���R��S{QY��7v�?t�ܰ����ֶJ������P�k����:j��`\��i+Kܚ0nd��?MA^h蓣8�v��<\�&���^�/ͨ�l}�A� lP�i�w���h	��Tal�%�wJ��˼��8��Cd̐��o�[��7n�O6�7��7���훤�Z��!
��j�7�@&���4���}g5����ᗳ��a��Y�00�����yI�	�}3����Ɵ'�
=\S!k˝9c�0I����]�[�G�i��8�����]Ct$��]�����/�;pλ^p-���%�����5�;aK�Y;�o��c��嗬}����i��֭�6��4����s��s��l�J��ZRL&S��Y�&4�ً��n�3�u��hp�a�р���KxKC^�)c�;����e��7thVFz-�W�e����b��ln�CI��7sMw`P����KK%��>��	�/b�I�Yww��#�%8��*#vrQ�H[��%��_��X��^���z@��Z���w9����@�@��\ǰ�X�/��	{��C)K�k�H���i�<�F�;��7�=�f�C[�T�@����3b\�Gv�I ��RL��Pl��Z�'l:2���-���Ntm�j���q�f�WsQ���eu`(��ڮ����Zy�x�E�N�R�y��I�8n����Ü�nQ�-�x��|��}�ޒ��uq�Y��Vi]�:���I�ϻA�$��)*�]��t�s�N������eͰ��u1���n��o�t^7��Ϲ���F�[�$;͓��C��;|$,v�"!wv� іk�;R����P5;sX���k:�]��cىuZu�йؖ�`�6�H�A�˨ި1	hI�hd=J!zp�un�}��$�����n��Z�[1��=�k�w�ݻ�u76���&�^�����۩vL\u�S��;Ӱq��zn�)*�Skb��ç����0�:nEA�g-��|�͢�i��ji�Й2�+}ؖ��;u`�Z{fږ�;������Z��hY�NM��Os�r���V��<w�DN��yn�\ku���m�v;��ʊ�8 -�&�1�˼c��4g\���n�T+;8��c�l<`��ټҺ?XuaN+�M������th���Å@�Ǽ0��pܰ;�sH���Ӯp���O*V��LΖ-ކSJx�W���v� g~�&"l�f��J�W�q��>�xp.�)�׍���<�3��G
Yٹ28wr�!�]����,e��\�it����oX�Y���|�]��>|s`Jw�3q����bozw.�����K}�."���T���4WZ9X4N#�h\�v�e>��V�q��"�4��x�d��ݑ^P����8wz�M����?v��˟� s/BΦ�*�f.�7��흽��:�̷tŦm��g)���fN�ׂ3��hB�>}_W��K'u\�|7m:���4u��cY���*SS �Ўpװ-Rd���k�m�S2�L;��oI�pt�܁�]Y�7�x.йc8m:�c��3��r"���y-ұ��]��zj�0nD9�?bk
��գ�z#@R-9H��NoH��o��!�^ㄮ��ٿ����y���c^۰�-�˭Y�ê���4H�~�}��ge��B>ٚ����hή�����ރh�3Gh甚�T�F\����6�]�tk�r���4�m���7�/ .:6<p��F�pi�1�C��n����!v�NR�
���dv�Hcw� ���K����r�A�݂q7t�J��Q�j��{�� ��ї�����Hl�,�qëJ�T���V���+���Þ�E}3�ÔQv�Cå�q�޻�>Qwc�j�&.��:�$�E�l8��c:�$z.�¶\L �e������˼V�šӽ����.���i��GE�y2f�$8D�����E�9*������0Oԝ���߄�oq�dT ������	^ە��@�U	p@�s��7���pY���Pz�v�?nt���@�kV^���c��-[R���>J����gM�cW6��_��ӱ��ʴ6�����1K�̺mcvk��۷�{x��zsg59Bv��LY*��@�6�
x־_��H���$���G!��׻n�w�j���؅lp�غj��������pC/C:� i[���f��v3vwvK�%�"Ŋ.�z���7CQc�7:dW:kV�Y����Tї�?�Gf����y����C����{^����D�E�p�N,=�T}\˖�+5���:����M]�P���Sn���Q��c���@W��cS�I��oR+�KC�ŀ����{��]4>���[Gn����3��a��:�wr7O~����:��,�,Ju��W��s{M������y���w�jt�O�ے/�W2Ι�+�Ƞ���s�%ב��2��}&����t��պ/\�ď�;�c׽+H��)��:*�7Y�&�TV��s�9ug0)%;X��;Z�3�	ɷAuc�<���ܚ���b�bVE�Ob�ӽm�������<#�k`�nx����CM���k���᡺�yc4�������k�f��;�`=zl+���0�Α�7r0��\���{z��$�W������+��81p�U�&Sױ���Y��E�=�ٳL�kWv�s{BZw\��n	\;{K�;7$�yLc(�WF�眆�Vno`�ѩd%�f�ˇo$�@���7�W��0^�8�/���ag9�w�T��.Ե0��T����8������7���);�[�Y.�;�9�V0��h��w���x,��E���{W �O�GvL�ܮ,����֙PKh0���v��M�+Mr��.Ń�@���vvFr�e��xMA�ݻ���GTo�{#s��l�	���X�1�÷�x�
��$�5���.�Nsn���*X#܇��Q�Û��Oo;���VJ�_�<�/��%�u�f6���̸���5�,RS�n�H�gq���:y׫��N�^�;�1wsw7M�{7z��@�����^α�s�j�{��p�q�q�՝��I�����ݷ6��wc2՗�Qq��&-k���KRc_�VΦr[y���SL��Ӑ<Vgn�VEO��`3�˃6��U-�)6ގ�suS�x,j�A��`���)��7��`:�]l�$�WH���i���|�,�F��S���;��T]{4��y�ב�qK�yn7�i��PL����a�Ԭ�x4�� ��m:�;��<Woty�0��UÄ�3V�gf�����n\�k��
Dx!�=3w�ʲR���=6�lgu�8���';�:�ݚ�sp`$�O�֎��;f�}�)E%�8C�S{f}�7(m���1��S���p��^��»��֖,Kۺz$V����+Ǜ;%��gt�C�n�U�M�=�p�����S��8�3@�C9�#g�{%�1m^5�.]�:�ҜӶoe�䚸��Ÿc)��or���F��12�=��O(o�O��oA�DV��ց� Kf��"���e��ټ�ɹS�HUw��p?�-�fr͹�iY1vt��lwV��,.^���-�B�����s,� �5�-w�.g��3�CM蹽چ��W6�7�-*�n��x���+^K��=�������}�n�I����e�W�������G�]���ܼ�l�V�8�,�`��3{��˸���b�q�Ȇ��c"�0-�Zރza�'dqΐ� (O�����9:�N�����0>a����u�q������N��h�nM�S7���9��.�r�	fS�8j�)q:�cǕ��D��[�p�;�X�_��=��0��6�Tn�ʚ���dU� r7r.�ýe�#��y��(�1zS
nڕ�'n�k�m�ǒ��������b�,��h����k�ޚ#U+�Ѻ��Zb�X�n4�>mɋ��u�s(qѸ��M���$���ȱWۯX����"#9z~4s3r�&�!�6�Xyt�1@F2�s���	��9�t���yđ���$}F�5u#�y�$t7�� r|�_�Ně=ӟh�qW��\O�ZNq�������؃�פ �PIv�n;�r4�#ٖ�N��C+�7��ns%~���)]���]��q��nѻ�)�)��ׄJ0�f��]B�ˡ����0���w&����|�ws�7N;8��0\sr.�v�\�����o��֎����P�?�[ur�K,��h�]��u~y�D�]2#�2�=��ם3q�*8x8l̮���sJ�wh{�H��p�ӻ	�r����s�ֵ��;���=\��{8���5I��1�,� X�Q)���`z�>���$seY,��p�A��.SA�ދ.ܼ�T�T���S@-�x���DѦiF��3WG��r��[�f[�Nq�̍?�]�X�;׫��X��eD��5�+�>F,N%7#���z�:��\����Ŷh�gqxgu�v��Tg.R��,n^�4�,#&=Y�Nw�)��aG�=;�Ԃ�ו�YJ�u�yg= ��0ê��7t�[�m͂�G�ۺ��W�A��;��=oj��f�P�G��FF�	��n˓8PY�,�hgR��f�?KIw5r���~8����I�^�oQz��9��X-Kkݑ�@����Y�$�q��\՗@c��:rd�j��ε$NqX��:�N��@�̞:<�ӯ9ۺ���4צf���خ\����2�BU��9 �C�M�2C�laN�w�]���!����+����{3r��������" ��:t~|�H�n<1;S��on=�y�*]{��G�kŸ�ʧ�ol���Ʀ �Q9j�E�����m����b�7�(���wl�y���n\xs����%��r�ǁ�{ =�ly^h,)Q���U�Yӭ��!��ҝ�auK��^�=��vcZ��<<ػ���4 H�긣7(�Q�O]0lf	�-��d't3ûb�V�*���[�Ļ��;#��KuZ��ŝUvLo�	S[��c��Wo�����v���J����{�7mK�&?�3K�$Nr�qE���ŉ]zJ$�c�q.��Ѽ�
5fMei�XΜOv==f�@�T���Gx"��d��MG�[�̻���6j���րV.B0�FI
�X�Cd-tΠug�Nu�×��d���q��/%ŏ8~X�����?�U��K�ek+���?�\��E,���r&��F�ô�o��x0Z�uu���}��&��_WǸQ��Er��{z����B����8#�&�������`�Pe]�;�Z�M\��$�ߞ¶lA���t��wJ�Y}��]f��7���-KI���#�q��D��ab�x��z,�a��
����L��v�?�q3�06��j�8��:����'$�YV]}l�ܴS}���b\G�h�(6h	7��a��u�0�{�^��nE�Lv��_�{�!���o]{�3�u"�n摝��[5�Лއ^���E�E*"��]��~t#I�sA@�mh�WI�rqO�7pD7h΁�b�r��u�C9J�VH&w��Ч
V�,U7�#�b�:V.��;L�\ ���mE2�iX��݇[�Ӎ�Fړ���u/ѡ����r�ˤ$0	�P΋x�Dt���r���^�%�;㋗"L1n�f�9dy�:b�E�4��d�s����2�:���T���)Q�.REY׀aDG_h��
+Cy�5pխ����V[9�`r���#΍��'n��o���twV��
�@v�$h*$��Sr󎫷���n�Y�����t���1���y�{�Z��"4k0Im]Ϣf�{9_:�M�wU���ѵ���Ν��ꍢ���d%c�wyr|_Ǩ��f�:`-�ez�r`�06����2���ÿ@n=����ti�߸�[�l#��b̔�f�s��.�۫s�;oq�y�RF�b�էK'p6ss�ٽ�Z�'�F�T�Q棗�Y�<Rm��H����:@�y�.�G,Z�N�$��9�)+��LL����S�iq��VR�^�oZeT��[<ܕ���3�v��K��׬�V�J��,Kyz-�?m�+�k�� �{C�ٔ3�^Ѻ���7��J��<�-��٠�`�;��d=R�^�2��9���b���ǳb%��7���	��lވ��r�V\_���L�L���Ͽp�e��W�CG�c?�?������q������?���'ox����<,���^�qXb���8�qؽ�0�-�-�%(�bib3Y)*� �V�u[1��p�᠔��t�.kƄd�D�x��l#,�"�+�ʺl�jh����^q�1ՙ�����B��tn"d�5�0���A-����Y`�Z[JU�T�ɭ�X��iltPð��qr*&tMu��(%�ɋj�w���W$��z�#69ƚbԙ� E���5c ,�J[��CFi)�[��du�)�l��{QYy4̤JP+Y�{@�{iTf̳U	BJ��Y[*B&�H�%o�4pl��y���k���	ak.��[���3bg\D�]�R鵶\��*�a�#eU6c,`ݡ!;d�	��ȨlJM�ƴ˅v�[��b쑦\FQ��˴J������W6�0e
P�3\�і31�dYSqix���WRi�m\qcҐ�<���dt�X�-���ʜ��qf�j����&M=�n�Ұ-�5S77��j0\Ueݲ����i���!^7a�ַJ��:6�:�F�j�i]0�3��$�[���Bm^
�J�ͮ�n��<���+M�������av1�T	[n�v�m�� h�J�4!t�S�'�8/��V�tK[h�J�J�/.%��.#H��髕�K�CYc0��3F�q6nX�,��5	n�����B4�\W3�U!���,�����pY��1����z�.X<m)�qYz��1�#T����Gfas���,�x�*�itu��BCB��]H1Xa-\��3�)I�5�u�a��n\P�	�S`*��-�lxf��K�.pS6�6f�݀ҐF�t�l�_�p����[n�"h�.+mQX�4WD��Zi�.�%n�;͘l(b˛��DM��J�4ʆ�4�XE��!Uݮ��Ȯ7^*��J3<f��ג�7���Pļ���Jܕi�kp�k�v��^cT��e�]R���ם��<��Gɻ��Q�ٻ.�4�q�u���PT9^�n���x�.��i����v�-+c[b;1�`ڸ��ks�è6�f�b��lC��k<���g��\U6����t��Jh]�v#1��f�q��!Pu!Z��l�]6ukl(�p.���t���s�U�5%�mr�]�-a�p�=mLf�	h��1sÚ8��K�Rj��-�,
��[-*+]��E��*�@�����z��Mk��P�K.̆�-����r�l�ƭA�Vmn�nD
hלa/i�؈˛ ��ZZ�,,��R�`������#�RR�%R;\��WJY����sjb5s�XJ�L���cG\�9�#��D�,՛�s*MK�pf�
�˳��.a�i��:�Jaɮ0���0�5,m�� �0ݰ��½l�S%�UbZ����Ͷ\�����1e�CV�������������]P�jƌ��ɭ��f�:k�5��$�X2si�[��b�A�[�/���ǝh�#Gh�b�?�����R<���ml)esI왖�RZ�&����A�g4�2�9�A������Sh�`�h�&�7�Ew.r��Yl���Q�Kv<���=/�[-mK��(T� VUIv��;���s�����D-�����n΍��r;X�Myf.0�3W��	���a���4��f�F(*dcm�( ��n.�Yr���0(;-�+	�t3K���2�2�h�5�ɖ��u�33@	��H3D	{��4�"�k�bl�YSM������d�(kذң����m�՛�U�:^��{�%Κ\�n�c0P�KC4��l�͛-�N.�2�sϟm��v�)�]Im�#�a�h.�ױj1��.5���i���2�7�6�-CYj �a.�l�+@�Ek�m(�L]�XRR0��<��d Km��\�'�	�h����x�J��T��,��D�lˈK*�0��n�]j�1#3����	,�ҖT�.6ɘ�b
�{舒1���$3��shEv��[.�	���5�ؚךݞ�nv#�We�6���"qq3�0qn띘�M�%&��m�5��@��L@(�\"�t\��mf"�L��YhZ@ԨE4�0�V�[bJ3]b5F.��\	��@n��G �-a��`�ܤ�9�����@ŋ2+u,��洕qV�ٔf�&����W�l�e�����6�$��V�4R"ˊ�5�����r��n�H�V���k*�(Dǽ���+�-�;i��q�Yz�Z��9��X�uxIZl�C4Ŏh��lF�1Nl���1���Ȁ�InkqU���n%�-�UC1�^f�Sf��u�5���0kd)�m��HE�8���Ŕ(Ǝ�+�F1�1i��l<�6�W&ejCsT�r�il
0����T�n�b�e�"�M,$W0�5��.n9�0�mC�,�sPZ�2�.GU�݃Wb��v{���K���M��%��B�#q�m�l���(���R���K�K��)	��菟hk�TZ�W[ҹ�f�\�V���;[*6�i�,���7�ڤ��L��,�Å&�ŌV��Mr�Q%�-Q�9KSiE��eJ6]Q�n]�Y�-ٿ<�=j�f��S"�#���݊"kQ�RhXV��G0�V�F�; �64���CY�-ج-MccY���ki�\b+4�	T2Gqe3zֲ�����i��i��T�6��B���\[�3.�1s���0�5����۫F땄�ņ�1BY�Ε&����3[0�[p�͛2%��#%3k5֩����0An��5��`l�l�Z5�
kG��C37&.�T��ٍ���"E����[�r���HF�fmŖH[.T�YuPn�m4F2M�M�
����mf ^V��cI�pF
�j�eJa&x���I�����B!E̓vff��鋱^���su"��� ;�me 26��QV|4_p64�6$ġ
�K%�7p�!�u-]5��Y"���8�slc�a��L�VXJKevP�KuּGQ���A���Z����f�]�����Y�n����"fXL��Ye٣nf:��k2ժ2��W��CUj�,3�v�)w,�iR,�4@��.j���ƙG,NїBU���n��kˠ��E�F����������v��HR�wЃ��nnl�K@���b��-!�l�%]��:����V�`�M�XYH�Xn�K�����5\��4��8��U��cJ��-�8��n���Vf&t˭�y2Xsj3J3uM��v���a�3-n��&m͆�u�Q
F,lR�d�h����#M��C].���3qG:�\�d#VP��#�mR�9�4��ͩ5�-R����� �us�5���xk���Lˠ䭘��c���z�g0ɢ-��[����@�Ɓ50ĳgb�CmY6�"@ֆ�����D��v&�Lv�n4c�h����K��S6�)�܄�t�Z��l������XqaD۞!,0�au
須��%n����6��;(Ϋ#(���GiF��L�m�5õ�ƁJ�j\ 9m���c�Ѵ]bi�)[��mEк�[��`K]-v�W�+iV��L�h��)�LfD Ў�*5��ԥj�W=�����Y��et%�g�,ķ���vuSU&��\۸��3��Dydbe\�WLL�X����qaq��+M�΄#3�Ivl��&�3M�DKÊ��L��hR%�.n��-#A)����e�F�2�ut#e�١���h���GL�ܖ����̑�1�e��ޫ�9qiQ�l�M	`M�[-շ�qqв�R�ն:��Z�PSCB8�.�XX�:ڂ�0��M��,�a�@�X�6l�[H9�䆹1��"�P�m�qM�� :5����i��5�8��
FlZgd�l�.�r
R+T��4YI���%���JŚS�iD���[3�y��3�e,�mu
�9�Mo^�
Lͪ��4�ג7k���� �]��e�������m-�6jí����g��ю����Z�I��6��,]���-�ih�f�f�*�W9%��B�]��MN��]H0�b�u�A6��z�D��aY5ˈ��Bg.2���f�Ry�6���GjhG#��ĺu�:c���.��c8o;fiB�b�!w+Y�������RS�"e��p��Rl4�,u-C;W �q� �جC)��8A,�%���Yc�(4T�zVVd,ݹt��v�er�X�� eݝ��Pnv�- �-� h%��Ei���t\!N�e�t@�\�f2���.�ք�2�����k\#\Pb��e�F����F5WL&Īi��2\�8���t��uL��FUҤZ�U�[�$�k
vcq)�˱դ�X/���C6� �6j bĶ:Lm�@F��qk#3y�*f�-�ڭ�#h��G�/7lW�4�۰WC�[�s�a�P�5Muk3��[X5��1r�Պ:��,a� ��V�B��2���6!,H�4��Dq��%�V��R�gJ�WL�r��A01����4-��F�]Yp���-�˙LI�)��`�����eY�Bb��Y���#�E�XKɪT��JS1ʺRh܆\��a��b8�v�i�*F�&��.���J�$U��--
�����^�Z�-�F696���l�\����ikH���*13�ĳ+-�kj�:�۶���MK-�3�D5�1KJ.�WV2�i��via�s�XR4��rMG��h&�Ή�60�e�kKe6#����[X�рj�Mȕl�[mx���mX���dx��\5�,�%&i�@��ʋ�Z����2Bn��,�DG�F���-]�u�n�S�ۇ��4�ѬH\P ����i!JϿ��w\^>�~�{���RU��������U���}��<���|���]�v��F�0���_����� �>�Ӡ^��Y����0B���h��M" +bl���XV��#ѱ0&�YXVm�X�d@z௠w����%���L�s���xa�O^��=����	��\�9�{ݲ=V����q@�J�{-K@�J��懝�+��,i'�Cv����A�/��p�6Ċ)�r��C�4y�|�L��}�<I�@F_˷7}<�{g�G���8Ԍ>h����"��ٻܩ�j��g��\��ι?�]��4�S������Q�}�`�01@��3����<��;�چ�z�)���R矏{�Y6����y�8}�<��ܛx�Kș��d�!:xu��簉Nj�ю5N�1xT�&�R��;Izyh����~�z�u����5��Qjڣ�`�L\�ȼ/nڻ)�#7��q�9��9Hd�O����u{{R�or������*�IW׺���}�Qrڷ��7��؎�?=�z�|�.97��_��{�1����^	r� f.�a�ڹ��ў�z�ٜ����>ۅE�g��=w�ڼs\�r�"�:Yf�d��-=gT,�0(�͂-z�T]6�r6���s,I��M��9�Y컹&�����+�7��.kʁ0��Ѱ�u�!�Tn�M���;�ɁO�<(D���<rb�P}w�.�*��O\��㠌��ͭG��G��o>��}�����;жE:�{�My��Y4(^��N��%D���53�!���g����RE�ű[�,�2�o�f*�q��x��O4w{���� GV'r���{¨�X��Vn��Z��1o�5T��4�8Bx����k�ߚ#˜[����~[�v��������c�^>�魽��`���۞�YW�YܳGn�x�ϳ[���k]/P�n^]@�7Fcc+a������������qj�v�7V#�}rxk��3:��j�gw/I�I�n�.[����;��L"껁(/���@yG��eػ'ˣ�*��ݸ��K��<X��t�;;�z���ab�s�_��8��f�`���Ƿݜ&��v��u��w}���_W�����~�x��{w7�<�2�KO/������1v	��?S�B{��2�?nrv�h�լ�艜]��/N!�w�T]�-��6ӄ�������x�z��FɧKcgC��ˡjC��b����������u�u?�f{�>[�/���T9�ejP�0��CQ3�"u�E��U��W��{�txVz��ǻ�S�PC#�̏H����6�寬~G�l�Xt`38@;��D'�WϨ����wz>r�=Ӯ�ݼX��ݗ�,��0Cq�K��q�M���9�cIu�5�W~s3�*HIX fR�����u�sn��{�^�!���E{��&_k{��]�]�͝۴dFm�І,ٽ��o�2�yj�V�������\��J�4�;��	4�Dm�;�j� ����wS�*�^"Z�f��z�D�ՠy���{�@�H'�8�;=�<q:8�"�/Wg�)�:3g���؇�˚���m������^m�%4���t���Xn]4՛�,�K�U{@�h^�]d�� Y��/�����m֒��z�؋cu\jԢ�<j�ᇱ�M���$-{��գ�ڲ�i�=����k?����Mr���9�����zi�E�h���<q�vޚ�����nvT�S6��V�/1Ͷ2��8i�.0�	 ��3*�N�m�L��^�P����j��w��!���.�Y��D�B�f���.���s�k�T/wuE�"&�g���O���Cħ4�N=�����W3o�	��A�:4��ϴ >;ey�i���⧫9��Oo,� fW�]�9��96�,��$�/b��|��D�`�_{��c*7��m�l�#;�ғ�Ym��se�Նc;��,YV���K.�!�.�c� �J�cuOm-C����ú�14B%@2M��M�>����AV�����|�/�b�_t���t�\��k�ڋ�J~�mb䮱����,[�^z�O�u��u�wP9v��[�a�@�"�h��~��P
+7:�� ���z��G��v����r�:ѥ��W���YF�J����a�,�k�
[Q"fL�hH.,M��a�5������W&�9�]�s�xrU��A�=S�40�מ�)��K/� ����Q��^��{)F�=|���D�[0���T��
�J�;U{Jvlc�����8)��"�K�&���r��ĸ����1����A�^o�s'���K��߼5MG�)җs��g�h�ح��r3J�J���2x<�΍@�PS���Ή�ﴦC��{R��=����	�%tk��θ�W�]b(f2�I��� ��y��\!$5�NN�W�6���yt_(��վ���K��v�Y;�߶
.s�l���[�M���������Y��������U�VK��6���AP¢n�v�&�Jv�R�茘h+(�b����M���~��T�����!������#.&�s�o�R��lQ�}��y��v�āT7C�4MFP��q�F�VI��Wy�icV���&P��8(�tm�O�K3ڗ7u̯�7�m�6���|q��u���kt]�ߓ��hzg���t$W��P�ñx�2�OD����. �_y$;��ڷa#U��}��&�"��,4�t�2R�`�+("��qT�����Z�lm�S��D����5�{��[\�����fƷ˭�����b��j$e^,1�L��O�tĔJV�21�a]e�Mnԉl㧫v�l<�M:uN���;�L��N�8����7�	�ۅ/'��q�^f���΍þ��!]Q�SNyoo�^kO��߰�v�x9��ĵ�]�.�]�E޾�Wbx�S��R�Ѳ|�J��y�(]�W^�/sc�˷� ~$��VJ�ۉb£ܫv��u�
���������7N�H���/��0H/>��a�w�����3�g�.L���0U�W� ˤs�~���f{�k��R���O�d[�>���_�r��~����n��'b��@�J�|=���f髓�.�O]��醄Oi�pL�9⣈<��Ch�S���q��w#GL�I|]�H���\��x�����~�V��S'|Jot��/���kթ�y���ܪ�{R�ӻA�o!b�U��ػ-T;�p�����K�cܤ'ӫ'x����Pb&�n{����e���_vv�R���8��u=��b�,҇h}�e�ѐ��ǋ�,���xh�$po�=��?2q~8�'��a�2BtM�A��7���zwg�]���a����?y��s��ժ�<[wH�c6^i{C1�NT-�db�5�b��}k��Ă@�����-�b�OF"p����:�I�D���0]�:ozu\��Y/�,����X��0��=���k��>~( �Qkg�/Og<F{_?^^�ۯQ���p�e�qBKwqJe�ހ�]A�H��:��F|��n����	v��~{5�i���1���.{4.8w	{�&�ێ��{���0���5IZbV	�qŦ@�<����QV@�9�2�\�/K�q;�Y+u��ǚҗO���u,`{��?l�XA�?����)���
���cu�w�:M�3w;�g����	#.�Nv4��|Y̙��z���*h�3�i���xƘ�!������5J쵲��3Q��ڜr�����7�̢U�v�T^K'���q���;�3/����{��}�B����m\�c(922Dlʽzg^��t���v��|����m}�^�oY�f࡮}�"����M���d�
q�90�ֹN���N�����X�hҮ%C�g���r����쏰�,�D$��~�z�n$�ډ��ћ�l��fm5�Fz�x���}t�w��39�è����ЧK�Ao���A>�"�SCo8qv5�+�=���^���#P��`�Z�ĭ��F�i�+"XWQ�k�Me2u\��jX��k�wuv)�T�3�G舊׮�[�=�y�w�Q�-�Y�Tܐ�F3"�[-���K����� }��w$��/RU�ŻW
Ї}�Y���]����@���*�Ot���;}�d��\�6bmܪ�y��0�)շX�XP�W%u��r��/v�p���F��|�Ob>:�r5��QRp)y�g�f��Lc���o���Zi��F������=�%xGv������ZZ���1�e��91��s��F�a�W��L_G�/}�C7�vO�N�FyI��'/y��Ms��s�;��9�B������i�+D�K���į��A
�N�\�Kܲ$R�b�p̷��D�����OXu2OL����8��ˆ���n���a�+w6e��=g�Ņ���Ӛ&%W��\��_#;Sռe�{`3	z�_h���>�5ǰ7�Z�a������ۄ+�we�ĕ�Dݞr�)���NkrD�ढ!��K���)x⬬³6�7�J	z��8���W/���fBF� x���l�ck7��t��4Í^� ��4�-��%Å2�ܓAԵ��"�|���ױb#��[�t-\��&�Aw
���ɞ��7{��g���^ʽ�	�[�@�.wX������z�'�F��|��^ig>�7Ǣyh@��{ q�\��ӧ��&{w��]��g�ص�w(�H8`��;�9e���Լӳ��a�Sڹ���{��f���������d\1Iȴ�ԝ�n������NK�8(AQSm��M=���c�0���q^U'���{Ͽ\\M�h������:w�͞�*��:{�/w�Y�a�Ƃ�7.���R���We��1�9�7i��H��ٞ���ty�o}j�N�O�ش�GV���'��{�:܊)�Çp
u��tm�$*�5��-0J��mM��5�Aٞ!���&����U�;��f)�;�@��é/cɞ�:���m�0���ӽ�SM��X�݃p�L9��~��h���b�z��r�ӫ���O>����k
�@��=6��սK|zL���j��-��oEG!U}��<BOg<��������~<�%Ǳٜ�E^&l'$e��k�h��cf�֜�fG;K��7�Da=c�边I������jj�Z��k^Հ�'�ƃ��j�6؈x]�T�ݩ*&v.�g��a5e�/���;YS��$���w�Q�O��ˌ^s��Fz��n���:���+ɟ#J�3뗌+����% ����t>9�F��V*�<}cL�����M�e�w.��w����=��%�+͞��''gR"7����w�g��1�=�i�Z{����{�8G�os ���or�o0�S ���
U��Bf�J{&��ڇ��#�y���]��gyc�%7̛�('rW_��#$����Fhar_Lk}�F7�2cJz�ۼN��i9O��x�mp#�Q��#UC/,�U5�ϧ-k1�ҳ�����k��w��M�=� �<�[�{�??p˚�{�<!����O��[�|}���h�Z����X��{ޡ4�iS�
��͍K�T[۹:�tI1��`X�*4^Xx�YY*�8���-���#�M��[����?6 ��w:��er�H��c�#���"���qP��օ���,"�|�k
��r�`��i��� B�����i۱o��gx��,�X��8D����u{��قip���{�t�>���,V�b{Z
��_�nE���漏b�׻�ܛ���dy`�zt_ q����=xL��[8
�C�|��ݶf	2`2Ѓ�Em����j�o�魎ק��C���B``��yx(a��:���Z��QƦ�<��(��sB� ���ge���I�RSk&�˦��X;�C�">֯�	��7�����/�����ƽ��Dxyc4�@�p��g��yӴ��gٳ)�67����N꘮��s5�0 �����}(�?)ȏ,j�С{u�z��k}A�G��5����O�`k�K�4��5j>��F�@Ϟl[��Y�}�p�.=;�.s����_f��Ѷ݌=[%z��jZW��N��Q������˼���k��3�G{�j�ym�;��1<��cN��Sxh��#�?Q�����.���t��gפ֕�Va�j�X3^�FP�-��4fq0Oma�V,� ��7����u�t��W���<>9on�=�N9��r�}��?�}5v��p�5�Ʈ�FA�Pw���!��y�o��_c��ڀ�뗜�ۯT��'��#�"Du��(ϳ[6�`}����1��C곸����tm[�[I�Ȫ,Vc�����ggh �g�oE5d���,Xo�S�u�{��S��SK=�=P��ӗ8�l��*�Z\1WW2�b�ۃ���뗂���p��}ܤ̂#�þ��,�-@�b��a��]&�YAV"�,��#1�t�R�}��N]���ٞz	���D:�fJCq���u�r�4�Vi��$#w%��|�Dj�_)0�ywC�\�@9g�`�D��D������1�˓Z~�e��{�Y�����9����w����)cѩa��4pH�Y[�a���i�3W����MIo�8�j����χ7�hn�}���{��3�L\bX�I�z�1o;��}f��]���;My��E��{&Y�z�Ѽ�sP�m��݇h~<B�>p,:�]�������w���@J�x'���0�E����Ә8�bMW�3Bá� ^��Q�y��<~���`�L�RD�5j�A�KeP�ؖj�@||;�ŜQ$�2����R�H�ޑ�;o���}�wg:[���|n�vs2{�ݷ8PWi,��K��@P�uqR���"��6v�m���h�Ün�*v'A4[��\�!a9}����+�t���yw���'�g�. �j��w�������g7�%wq�ܒsܛv��~�L���g�w��d�{`a(��Es��_d$Y���\p��=��w���]�u��u����=�}�Z�U�k{ni��1Ff�\�q��ѷ���T��lp��ع̫��{��6@D��0aYJ�h;����Sy[���Zb�t�;������+�d8�X�A>��2�n��5c��\"���w��$y�XZ���s�&-�uk���l\�܇�}PP�����k�L�..��?.�P�=��z�K(���?��>�EUikl������ݜ��|}o����z"�*������Xf��!	��2AD�6�Z*�TP�9�KM�zt�]6�ۅo��%�eݟ���?]S��ٙ�H|�Uĝw᯿��:��[8����ɛ��63�#����T΁�7�UD���o�ϲ�X����KI�xsZ)�E,Is
���ĭ��v��Z-�mX)l0�!FX����a v�ۙ��5���M.�ˢ�uQ.��@���ض�,l�i�1bܑkXEL�.�`�J�Zqj̉���h4�ƣG$f�`H�	��)s��-,K��@K��uB8�ca\�\`r�3��7	3h�L���x�[*��.�Wav�ۨ�b�����ٴThCl%5��3M��f��+bC���aXs�f�N1���#M�5�u�Za1�h�Y[U#,����7N������$�j���Vn�n�.��)�ةT�M+[����n lĐ�N*[bq5m�l�b���($�G*�kN�ն��J����Ȱ�ͭ�sV���c�Ȓ�d�\���(U�����i�2�1�T�ȱ�56�1Iv4�ƈ[TF˱�69K�����hB�1�2\Sl�F˙D���h��,MQn�FJ�,It��ֲ�MsT�s�!e��+��iL��V%�1����׮���h;ha-	� �Y��p즤ʹ,#,I(V�u*�]%�	��i����tD5�!�u8��̲�e���6��X�]P�)x��֑v�]q4%�"F�^�!m"j���ɉ�̓A�顰�ѭÒ��-@�żK��l�j�if�Б!@��k3Ҧ�k��-D��鮉�Y�ѮxB���aP��֠���<����Zͣ���KFlh�͙A��CM�a��$�0��15�NF5�cSJjq���$J�D�����]���kك�n՗�:�J%�)[LVָ���d7cF]����T":�PJCn����j��&��B�ä6,f�77 �2��J�i�]Z<�m���${s.ڮ���(£k���Į�K��%���HE�.�:�Iu�Q�#��jl 3ڷs,�YD��XΉ�a1�9J͙Jر2�bj)@�a1�B�oV�Ji�k;6�d�+�zEor���DK?�� vq�������5��S��g�873��U�pU7F����X��4\�4��o��rz����܍b�CGљ���_ڤ�A�[���1��7A������-<��]񮗢{���/���.无��>�z����N��ъ�A�6�fٰ���:{��[��d�#L�gE|c��&ll��p�/#L���w��<>���V1v�����o��u�ڸQT��E�����#��{�Q�/p��0;���(��&�;���FY�#Th
�jP�=^X��Ǯ4-�_�n��N65�&�"���c�k<n����&3�v��:�Y�{3�	˓jG_�j��2��1b�!�;s�ŗ�;K���F�c��Y�Z#d����>1��*_�O�|3�Q�_B�js�s:h܍L���񅛬M��B�V��f7ُN�D��=���d�j���\����9l�х�00�A�@���s��G�U��Ȏ��Z��>�dRZ�f�S����Q����wU]��o�x�v9�A�f�Իl]gVF��M	q���lr�$Xj;�U��'˰��+y��9�B5�G�p� r��u�`�.��������g{ln:��A[��/}9Ш,��ڻS�)����.U���	�8�/��/7"n\�Y�}�.m�f~Ѝ<���.�_����67tZ�qY�:Gzb���(�N��T蘽��j�@?m��߽�����3>��0&��T�m4M�x |*�E��<�sr(Nt!��{7LΙWx����z�끴:%=��N�գw�{.����������G��������t� Jv���X�(�i�SZ�2�J���lb1M��iYk���V6d4�!sl���V��1�J�� J���� �6�mq���2��8��S�ggKx�e�l�8��dv�l%�afwB�o`��!��t�,V�JJ��ƨ�h�0��ICM6��\�\&W�f4�̣u����	BB.D|�ͯvR�7�b�a�K�'͎a/C��ʹ#����z،���#��Ã4Q�f{e����6�����ĳD*�A��	ThDJ�U[5�N�1�J{���X	D�iϳ�.�>�?s�̧n���z����9�ٮ����s&bL�J�n�v{�����bAB�&�r����R�km�u/����� ��I���/�#���^�î���'��u-�����bK�- �B)I0�u�/�ᤏy�3k��)5�\�e�m� P{��	����%�L8� �m��ya<x���{|6{������22�e���Q�o��h��.f��++eBksR��7I��%U��o:�.
�`t�3f���k؎ʦ�m-h���l��9"����{�=gâ8�qpԽ\��>0��
H��p��+5�ܵ9�-S�o"K3n&�q�ƀ��Q�!�$�Uz�;g�8d�v��8i�[}�t��žnۣQd���%����QBU1�綒�P�U����vI�G�̺R�dA�`�K�d#oz�YT��*��ƀחQn-��Za�jT�
n�0���-��az�b
��`�����S��J;���>̴ӛv�u8��u�	%" �&"%+���y��{-Lc�x��ʍ��vp��Dy��p��5dp�&�L��N#��ѳ�zG��W�v\��Vm�ˠ����~�p��1&G${&�v��-˗0���w2$7YJ�E��5���|l��Z	��-68Ϝ��3k�;'N��_���8�Lc��B��&@�D̔
Hmmdk����3�5k�b�&/��;��1O�@�`}�H��)��\�Og+�{�gw��V�P�1�vE�Ț�{����{�lt輄1��7	}��C|��v�x�g]H�ۓ��tի~W}:y�Q�z��;?l�,���~�_0^P�3����5G�6�|�m�\&e~�Wy{R��Ƀ���9=�쯄~�	0[$�cqz!`k?~�3�t��o���E狃6&B��H)$5w��[M�<M_U��ܭ�Mn8�g '���}=i�D�+�d�����;��������v:�Z"��ҋ�+V]g{�Y#&a�ƳJّ�.�Ŧ����n9Bkr�:�u����l�D�I��Wj��ٲ����}��x���&6u����_UOV�p��L	�&�$���R��؞���=n��s���N-�Nt�����"���1��;S��;f��@=�_����==<��>Έ��P+�`���C���|=��{%��x;2�W34�Ž�E�۫|,�w/c����3T���bE�b�<�1[y|��������U�rt��o�nľ[\)
�u[�=�鸷�β�W%��}?��Uw�R��vO�cDd���FA�ҙ�YZ�C�Xia�?6�{��K�8�������OC����� $d��R�R�h[�qp��z��-��i�F���uVWxxw`�1"U��̕��If�b(��jB��s`��J�+���jh�S$�*��UT�_��2�g�6��F�q-�<����U�9�`��fPI��kN3w��g��ע�W�rP�X��Χ��xW:y�M	��`�% �!��]pЭ���c��c�f�N9��7Ͼ\���9� ����%2�;��'�|)�솲���FU,ݹ��=��j_dUV��[$D��a)ӑ�������&5ˤ�8!F����=��/�Б/f!����8�:+eQEb��&c\m]���Y�Q"h��J1Mp�:f�s�C�t�h��,�;�v��+��{2�ϑb3z6�e��5�0A�:������cYiM�세��LFU�d�A�Yc�=R��;]ڔ�� Gfc���0k�7\��^e��gh����.�Y-Η��1Ք�+A����P�u*��]RB�\�s��7y��>6l�C:吋4)Y�[��1x��BՈktH�P��w9���e���M,j��P��ơu�ȑ��&��A�&��%�Vn�����?�PF��)�8������0�ָV��feʊ���!9�!
1�vv���������ăCG!��ɫ�Kl���P�ˈ�l�I�Ƶ�iD�e���8��@�e����~��w�ֹ׫=?��^�յ�I��X�	R2�T��P��������Ks[�X�A�Fl%s�������3��RJI�%BP�Q����z+d�댞� �z��Ơk֢F	���̉�>0�D�$3f;����46���×��:��l`�l�Д���������Q��އ;4{���_Om6����qR1b�����H�'�԰q�0kmf2cCb[�H�f�-ak��se/l�
XD,N���B�ޘ��2Ү���!���Y�ۭ��K���ު>�����fk�*#*T�JQ���z�2�5�Px��&n�ΔI�=bi
��Ċ���"}�"F�� "Q��:�����A�|���{�Fz�i��`�4����s$���8nHL$P��Aq ���d7�%?&�����{����!�������5ڸ��[��,0��":�\������Kxz|=[�&K�fH�1&L*�-eWST�7����������k�t�J(G������� �z�_d�vn*��;;:ڽ�����,�^�{h��H�fb@�%#�������G�r��|Z᳒ozk����������$V"nI[��Pn��a�q� �j\4�fփ,�V���,6l��N���Ӹ��ٱe��w�!�y�~�)}|��ˇ*�)*��2�Z##C� /xS{o��8_KN/&*s]*������l���
	J`I�1*���91�V�t0=y4�&5����k�%�b�t�tVle�/�IfwUR��S"v�#�H2ғ�/�	ݮ�}��>ᬍ�3#��â�R�^���C�D���1(��JgbjGy���݈h,,�������![m�ճ�^g����bc���̽��-�ꚥ�!"%%��w���]�Q�/��̼ة�֌������|}�"��g~�)��"�;!���1}�	�>F�+�scl��L�>}�M��;%јpV�m���b]L���Ը�
-�ͭ��]��.��ΟD	??O�},<@L���-��۪[�K-Է���Q������w�I� �&D�T�6p&���$����&��F��⽵�U� H��s�=$�T��锏S5<�ǣ(� ��c�LÓ�mZۧ6v����NS�ɉ�sG_>ȅȉ��x�Vt�����;��C*��E���eLU�)�@�.2��*���i�����d?��=��:s`'��a�.Y5��f3���\xI]�F*�o��qkףa�6j����N�1�F6��k�b$�Q�D�/��7��Ikc�u��Ћ+7V�A�$�s�<3?���q�^�e��a��q��::�o�����{��Ee��ϛ�1$���yХ8�-�T̹f1Tvu��4�����f�퍈���A��76A�,z"e&RC�y�};R�ь���q��s�_^x<�Z��~x�)��2�]�:SG4�{���b-����Ҍ���q�<�-��{*J!(��%i�k��ã����7-��o�;��(eb�DKe f")��7���}qX���K|��ËS�����=�]ӱ<���R*J�1338��Nwn������k����pnHW_�>�خ}D؇D�n��1�ux��Q��x�^�>\j�� �+���܀���� ��9I$a�� >�����6yK�Y��ٷ���=�������d<~ǀ�m C�a�����Rc��7m�l��4�
�/]����7�f�(�b��ұ�(�#2X���_۝��ꑇ��[��a[wf��a�P[/&e�ݵy�l�o0���qi	A���Y\Q[��%��i�^���C��]bͦjh���056�&�a"bS����j�٘T�\�R�Z�].�E,|�mڴ,�s�dş�� F���Z���H��m�g�ŻG�K�w��oKɫv���s���KО<�/��V�g���Z�X�H��kGTơKl��a�Yf����Z>,!t�����'��i��uM�}g��=qՃNh�d��J�*Zf�'ZY�=���%����\��f��N]Dw�� #E��Ͻ�|ID&_�l�>�1GZ��.��9=ˣ��C��w�Cp"."�AJB�L�Q�+�#�Re�����'w�vSd�GzG�ݖ6qh�:��R%L)
T$��j�6�+��G��ͩ��4�T���~?�z~Ο~{�~긙�0p��1ö�̛Bb=�M3�sjB��#^�A�K�2R�&�XS0�)I�T�}./����j_{�]"���-lj�#�bPE�*S���ޚJ�}�ZVWq8j����ё�[�7�)�p�����o�s���ju�s��}Ovg�E�t��2r,�T���fr��"�8D�sܝ��{�6pl~rvR�ij�S���f�Qm����!�n�"����{jB��ߘ~&�A��n�������u����62��997:��������N�b8&�e��m`I�Ӯ{��{7׊�;���~������;)���WY3"DIP�D��Q�;����v�κ=<�cF��x;������(f|vf8H���)�I���<�7�O���QQQ��՗���r{x�_�\d�bp1�	LsNd�9�ZFb�Kt�[�\�qv��j1Vi��Ґ���S	��)�OBᓋv]�Z�٦;����6v/��a\��8lM��8q~D��ź����  q����э���Ӯ��y���g�}����h�B`$�S�ɉl✼v�U�Y[��ɐ퉓sq;B��R�R�V����B�b��=��{ܩ�Z��>�wfz� [����,���o�J7������"m��Cݽ[G��to����'7-�^2��G���}FS�NI�[g���������}��䍻no�Y�F���ý�?%@����A��Cw�{�@x��Y�co�J-��{�%�TDA��4gd�x�|��q5v�X��R����H׶o7�����=<y/>k+U����Cj�{�fS�&��fcB�>�E�қQ��߈�͑���J5��c*���SV�ק"q�"J���]Ef��^��]D������g��|Q�V��<� O&	��د0E*���#0U�M��'��^�F3����8�Z=�~��_}7��$Z��T�e�u�Έ&]�$h�+��`��J,��ف�\Ԩ@r�F���;¢ީ	Ӽ�_E�G���&�*�"���/x/�d8��r; ���nKr��2l��)�����Q�)�?Q�G�ݬgx�Ȇ�� �OW�|�|�ln��ǂ��4&�e��m�L�J.�l+1WKIɻ���f��4�M���.yt��]��^�H�7�F����Qe�s˶j�la�*�2�)�|7l��0AY8K��QQf'���g:�F^�h9�Y˻���uO�e]N��g*�\DG>�7�b	�W��ڞ԰u���i=G�c�{^On
�LN�=T��7<�^�sھ�]Y�'o�y�Ȏ�3n]�z��}9b�YNo�����D1���#�/�O{nH���ƕ�rB��ݚ�B��
�%
���.���v��n��dK�G��ttX��Q�s���9ȕk!�1:x�-�0��U����[��up��gOQkR�=�ݷ��}�G���ٹ[����dj�����O�o �?�Q�y�J��4>���Az��޹����v'�es��:�ԧde�t���;�oH۾<p��vQ�k:�ਝZ:ع�����o=Irf� (fR�Jk�.0Fd.u~��x��n�뵀�l��Dg>i3#/�o��}wۛ������f�76i��6�8�P/k7�=YZi��k�]��|)=ӑ�*����K6��޶5���٩b�$;c.�E�S[�tW]k	
�v��D^)��X��Dk�=�u�b�|1�9ў���ѧE�42|�ֹsH�ֆv�Y�2vO�*��F��b)𚎎=�4z��{oR���b������h]��{�Y���S����.-g�G'ʳ�eh���kl͍//���TU��ow�^.9�-�ac��J,+�z,.)B]cׅ���4·��V%�U��M���%�o���;�z�g;"Ob&����fX>�~��N%Mჳ�j��VR���VH�o&w����_fN�����v��ewȯ�7���^3Z�}�δ>w�6oL�l�^���7ˌ���d�^01�'�"C�!lU�&��W��}]��_�˨0#e�4)��)n����M� �[��P��������#;^n�`������s��]�k/�51*`缆�k*��ڪ2#|2kz�zt>�,Pͪߐ9Ü�Ă�4�"���S���V�v�n��Ǧ̷f�?�I��"�8Q���=�(7w{�O�-��*tEƬ��.��w�)�ȼ؍�53o���������7v/fV�Cv	���؜4gH������
��C��{�:�c���8�����_t����՛�9=J��dD��Z��s1�������4mġ<S���&�0>9r�����K�!>4Ȉ��e���+<RIxP���*�V�ԛ�i�nnn���I�����TE�/�D%���u|0u����]����:�y�4�z��=K֓������;����=S֗[b��/�8�SN��Z�������b�Q�~;�y��{�믅u���y����ZI�)�P�s���)"D�����v�x�V/�aB��Ne��%K�*�4�&�n�B��b����TT홝.�`ֺ�>��=�����;W�?D��~N��N}�ɿ
</��g3J:D���Q��Ο	x��|7Z�rwχ~�|y:��>�E��A��6�
�>� �Q�	+��U�^��V���F�����i��<��p�E�ocW֢0XD.���n#�5B��Ia�fj��s%"�t�۩۞�u���{��W�}w�z��^sǞJI�{괣�M�P�'����w
4RD%�K��ۏ�
�"��cmL򩍒�2��]��q�\=��B���	��)��@���>�<*_8�4��� zgs�D`����-Iu\�y�Y�럾;��;�=��1.�4�DiBLӗQ[��w�y�>�숭�ROMB��I�m9=���x������t һ%����2���iȰ�Iݖ�>G�����a�&�����6`��������Pv�&�팄$��[�������G̏~xAU��]!/�de�l�C�NJw�zݼ�|���v��vz��W�8u��;�iԖw�P�	!.%��W	|+��޲�GN�|$�-؄��~���6R�����
Kf��B��0��.G6��[�K�ey�]�|�,jj&J�%7ussƒ𙂅B����n�h�O9�S�>��G��G�v��緾�Z�\�MG�KI.w��F�)u�_������fG%���Q"���%3�����%U�"I�ad��Q�(]#������-<$�
#��{�X,Ԓ�Q*8a"�����)���U7����#�7d%�o9��D.BVB^�x��EFwa.$�����Q�E{Y�Ҏ�$�I��E�10��R�Z���w�#�J�uDzZ��Fsw&�"!aD>��i.�ģ�I��T`�
"<.��Jb�]�9ڸK�QG�֓�H�PM1U�uwn�/	.q��T�;=�s��	x���]�"⧾����a��^�"���1�� ShG���dBF��{^����7�}7|�}יfnz@�zG*���3s d�(N\_VͰ��6c����ǝF)ڬ$����Ʒ��J�IIW�<.��2�Eh�B�_�����ff��r�*+rXfSE�;�4�ل:  �2̹��v(�j���T��ńs�T�b\�PI�������2�F8�a�Ku��<م
���JYD��
6�y �Y�����H�7^�	���֛��i�LZ�Xdti������"[��ް7�5BlhŇj!HȱȘq5�V�X��6I�M�]nAY[�,�H��}����������UFAq���'NNǿQ���nE&^�̚$��뾸o���M�m(��R��@�qaG$����w75;�!�t�4�h�y�m���6n0�hı3.5�YZo֞�{�%�.��&�����_}D��c׿����w�1�w��o}�C�s�GXz��ӳ��x\���s�Z�w�}��X��H���ѺO(s2ۙ�3p��Yk�K�}iGrr�Y�"�S𗄾���j�Q�2�q���	|G2�5�x{ �,�g������#s5B����ڼX�P�e{��0J�|섫/.mDN�%*%/�'J~�v��Y޵&niGE�%ä.�lN%2JJ�� E*����| #��dD��B�5�w7�\Y&G�d,���it�O�ԬH��GE��MF
$K'���?R�E"�һ���Ƽ�n/^~��������ڼ�v�|Qӂ���p�����,������&��p���\6"'ٳ+�[bmȦU�iX�sB�ȳ-.��[
!k��p�3EW�,�n�M�$�'�w�][c��s��~���:x�>�5�U��K��s��qH�(�5���ٴ��"�֗.ٚ�%�%G�K��ƜUT�r����7rr�.���1��k��k�s���)Oثl�=��b{s��7rIO��y�iU�QC�%�0P.�feU�25Ga�ѝY+�P Ix�T]�h���3���}�L�����6['��FPcr'<��k	ڱ�Jzk}�H'1I�=o���\^��U�6A�C߃���#�%�h�>dQ��#HݗCò����F֪�f������B�Y�1.|&8jS����!H��#�d�%b�#±,�{�7���Qi)�n!{v���/�R(�g5�G��E����%r�4ꤪ��wv�`�%�uB���"��mF
$��X�v��ixVYb^�n;��/�����S�ٵ"�
,�b����	���f�n0J���t�DZ|.��سb"R\����M���P�}���aB��9̴��#�E���Q�ǽj];��e�rm�K�(;�V��б��2�Ҏ���tEA�w~GXOi|�.��w�����I �(��t�>G��>	��x i��;�Z�Q�T)L���N#۵�-8s_ڨ.��T:�*�nݯ�KF|�|�W��J�}���O��NS���ԯ� Ȭ����G��c�(�諛��U1$���l�uun�)<���Ns���*���q�!�J��?�L�����D��%X�&:��EǙQ�]�꾨�:T�����d}u�8A�w[J�
������	X��/��p�`�}�����_k�)i�Ս�v�_�%9Y��"�
]�^������<�d��O�jV�W��,�����]~��ߎ��0�����|(�#2��3 �L�0��P*�W� 	1��⋅�C����K�G-ǻ�M(�ĺX�|W=6����@D)q�|ssz�.�O^��BJx�e��ne�7v��:�pI9�1߈K���T.D|D�>�O_9I�*8'~�^ $�u�8.�s�ix�"�J=�ٖ�P�D����Ci�)�t�2�83u#\JJF)ٸ�=T��<t7y��.���jݭ!QB�=ݩ�%"K���w�s}<a�r�E<�Q+���/��ߝ���DφqP5Njj��\ݫ�H���Y�g-,^؏�tR-S��h��>�P�"����y5�A��T�!*��O����F��%Sqnjˌ(]!1wr��a�GH���g�����RQe�u�~���t�
��I2<���(tI(����
g�}�$����ޑ"�p~��n��Y	ξ���D3���u�j#7�w�!f9M���ם��{k*���U���U���V����TI.�Oh<��#)�{YU�[9�h;�;)v�.\�d�VZ���3n�u��'�>\p�.�4OяZ^djRI�����i��k���A�������'E��`� ����^����I0�C�Q�q�&ce
����I���ǈ]"(Q9^�x(�;M|~%(�Kv��"�BU�y6�)$�}�q�D	X�E-�
p^��*f�n���Vc�4�L0��YaA-�a�R��d-̠҄Jm���;U�-hl����'����Է���p����Vrݯ���	��{��b1CA�����y�/ځ�)���m���4��t/�%�����؉�GyQ�{y�\t�	i��>�Q"]<X����,+R�IO͂�i�h�]:�D����Mia���Ϸ�q��G��*��q�sp{�%+�=pM�p���O� ϯU������`��qjd۪�X)Df^�MEGN�9��\FF.��)�/2<Da�n��L�(�E����7�J;�Zr�vH)9T��]��+��3��J^�Ӄ���O٦�-���mnM�λ��u���>�*��<&O}U#��醴�ܺ���D��j��Y�u\�Cw;%p�v"H×���)rH��K� �����4f��k�w�����&C!�52�F���	�!�V�Tk�;�bY)i\��K"Eۅ�ԉ�tƛ=�j�rM�2��i��1m�b,�X��љ��(2���[��m2]�@� h�-��u�	��Rf���ⷨ)mlf�b�#J�͚��[���wy<�{� ��L��,���n����z\꜑��Q�vAԬ�oX��t�ҫ�=��L�?h�gC\�-��WGN�H��ӻfwA_5�����c�����;�&&�^�[��F6�iX��Yvj�6�eK4�S���<��1�"E�kaE���5o�<|��ZmKT���	� p�S2p�>�בL�f����W��G��E�(�V^�0��Ф^������4�UU^GH������u�g����T�&,8G'}�|�)�2o�k�W	�`�����B)H2i����ջ�b}��X���g��q���
:�ş	L�1_��%fV{]���r���0����o&4�S1�~ g��4��U��>�����*H}�w�G����+۪ش�<|=��iUINi��J���a�(�g/*�RDZ�)X�{>ɻ^(Kォ�azD���ɼ��
O���^�}��IN��l8t�H�"mKu�F�H&���.5���f�M��d��]4�9U9uR)n��.#Fp]����p�Vp��Y,���-�������˘�dS4`���r%L��D��)(�>���}[����ko��f�l}����C�f/	�y�&7��Q�}o�(�S����γVt�2\[�Z��swF6wsS�u't�+Y�*z��g=������M������m��Y���߂�h�M��]� CM=�N���M������$;��E��[�/(�� �Dw6(q��A 4ԦQB�S����^�)�)a�<t1;z��JdS"sT����\��ǆx�=���U����',Zf�f�ā�|\��j���WqI!)EJ�I�-w��J�F�~�/N�n�97�8N�xGo׎���R��;��fx
ŞG�.�Ln�)U�_J �sry�E؈����W
��Y���q���7�A��ׇOl(W/�6�:l���)&�[-c<	4�ƁA��٥kf�����Aṥ�N��u��)�T�.i��O�b+n�sDt¸�]{HeP0�Î�U�� � Q�&�
E���y�N*�r��;I����}=��������[���wo�	x����}�+��O�3���K+ H,s�T��0A��:1;��J('�CO�+�d�<����얊�;:�^yܿ�����g�bY$9���!r�k�*1�Wl��"��
�RBxNN��#."m������9���h��>h�>xW��o7:w"�1-;<�䀡���rJnq�gLx�9@y�;���p]͚� `/�{�q��,�l��GTN�4Y��1ދ�!��]T��t؈�$��fo��Z�Qݫ�x.
�ز�9ix��/T/(�O9ݛ������7�޶�P��K�|*���3��b�Fsa/�\�ݞɥ�c�[����.̿��B�A����z,�9�y�hY�v�if��9�4*rY��-��`�.&NƜd6�����7�_>^��Yw_/Y����y�,�Gi��]��p�����ݿ��Q�Q��j�ʦܦL�sNiZ�x�K/*k/R�BW
���Ӝ:�a���p���L������ͅP��¬_���KT�Q.i^D*v�5�I,�{�v!)�ITE,:;��v,-	tK�����8.�X"Q�(���j��B���bqtἝ�~"�,���GK:���+�~8%�Gݬ}�4zr�eN���ɯ���uzا"HA�b ��'�w�oѸ6bC�3vY^X�T@���´��g���׍�9�$^dy�<�:�4�)���[4�S�X�w.6�����8�Og=��x۫P�[����`���PK?<K
�]U�b�!���S�h3dS�����A�2�l%���( o��Z��#'R��/����м/�����K'לW���	Ԓ�g�u9Mf  !JX�-���B.(�7V�T�!�gb99�f�R[7|8�*��.d��s5��&-��;��B�޿:�#:Y3�x��M$Ҝk�3y6����z�{I�#r��ʛ�un�\:.�g&׋�R"Tf>7�_�P4���װ��6D�6+Np��"2<tig����*duE+���zpX{菺�P�GL���������+:(�@�cn�-��@q򘀊����xaa�l@�m�s�߮4���zy�ح2|M�·�3��}�&�s@!�c|3�?�E$	- 2$r�
��q{�����_�=/�P��2+J7p0��^H��(�(���cq�f���c��n2�܋E�����(�W:�<�na*��Ӻ|��1P��	���Vm����\T�E��7��/1�gz8�잲*��J��kػ��Ԇ3tD\�A�J�,i��~��'dd�g�fp��wEW\���u�*��F	�<����C�q�\V_i7=�?+�C{Ǳ%�wl+A5Us���@��7A.E	����`βgM13s53�J8NVǲʪA�t7�x"D\�=�+/��U&'�4mgL�th��B�e�W�t�{�.m�U>���D+�ݭ�xz'^�K�Gw�p'=dw݋Ͽh���wRL�L���$	�[������]����g����'E�ċ.}��̞�f�=Ǫm��窛���81?s��$A������'>6�8�f���g����Ê�Z�W�.��.ڷs߷)]�	�u 6��Y�q�/�ٴ�w>,B�~���l83�<Oi�Q�;�n��9�m+��QJ�̋�ز?!�YG�������%F�I�	����c���'��0�����ꭓ�3K��L��mW8�_z�Q홋�+#��v\5�&�
�	��:��Jj�E+��^����+�:����xs��d����'�S����� ��u[Ӿ�
~��r�2۵7����FŬ�pC�1��_k;���r.>H���ML�ϗaL�aY����tn�\�|	�S�\�][<�ΰe+�0���wI�r�|.oT���uq�n�=
vMR�%�o����{/�W�INx��%E����e���Nﻼe�O��dj4b9��5e���h��r�~��\Y�Gx�5zd��#�^�U�tMC̪��j���T�wc�Vwf�r&/{h૖�U��q�7Ѩ�I�0OuWY�ȫ*e���^���R��`ʵ7ۨ�z6����&~ލ��0�.�K��ݵZ3E4�uc\\��f�i�1ٶ�	���C��ųhU�-݋�bf.v��
��f�ٜ\69�1��0�sٝF���s�hjk6Rۖ�iuCDma4hPc��:�[Eq���c:I����A��SWZG.���B3\�Y���݉���ڱ�Q-l��'V���v)dT����6z.6��v���Z-K��q�`m5�A�K�mMBh
�F�LֶZCd¦CBm����jJ޲�L��x�p:*��k���l�����16d[([#2�W8�m,/\�ˆ���ųF(�)i�\]+\�Vݘ��\u3�8�dD��M����c����.射��H��6au2Xcc�Kf�Ά
�C��7MN�Ս�,��bS ��2L�-��25���R��X�gvZD���{�ˠ
��F�	��Y��qB̚�j�JU�v�\����� `]�����������x\j�z�7ZMe�\�n:m
Ai-!��W5��h*���ຂ��C@�ʪ�kT5f�2�����č��f\�!�,����bWo2��O0"ͮH k3.qՅ���@B-2�Sp;��>i�|T4Z�ɚ;[JM�[B��g:��ûc�va�ю��K\�Lb�L�y��TA���q����wk�#uu�ѤZ!K�lR:cX@6�����Jg-��p�c͖��M�R�rB����kl��c�Lg����,�1���,ڡ	X��jՄ��IsT���f���N,M`̳m�R�ȓ0ld-v��M*��l-���`��ia�Y@P�`k�r��  =t�-��m�6��&��ad4�Ql�"�u�5ִ�h�����hG�k������wid�L�	�3)Q�.���#S7P���rk��A�e�IH�n�f;)cq�J`s�E�����2Lf[�Uv�4�ν�0jB� �Z�iYp�RfT�B}&f/� 3J�w��sm�X�?ng�a�O`S�ӹ��BҞޫ�k!����n&e(^
���M�FGep�w�:d��2A�5��s}��k���˞Ur*�և\�Wlm�s�G-w�7������&v�OS�����r�y@T�Vӓ�8,�����3��b�4�)s�t/M�+:�(����3ݢ�/���Ϫ�p�lj��!�ފZ&�
��ܧ2��X���b�N&{�Oe�u�A
��-��q۸�GarJK��0��'&d@�w�Jñ�r�Q:��(X0�p�E��M]���~�I�F�bE���r�48g�Ͼ�{��/,�LZ�ڮ�NC�F)�n���ǫD��oDފ�tE_���pS���9`Tɳ7yx*�#���O��s6�Ȉu*��Ms��$o�֩����T�|��Gqغ�u�ӝ�9vs�軝q��;Dc�������=t_#�v)���6kU8ֺzo�!m�֜�Q��kn�]��ͨda���~|V8�洞��� �T�$��s���=�&
����Sn�G���(.��s�y�&ı 5ul+�D�\h�D/�1yU��NG(�3��}af ă����{Q��t��*���L�3*T�\ta�Ż�8s+�U�؀�.�b�F�#8�j�%W+saZOg�1mN�a�t:{�p���L����
��{=�¨��-�(�U'NZ��������ʶ3��lύ�o������i��|�מ�W4v#9>��^�D+r P��[�L�3���]�q�q��lvQ�=�E��N���)�ףO�~+=9F��sZ�f��khU#X�R�jڣQ�\�����H�%�Kَٮ�6�%¨H6T��.���?�V'`��4ѺR��e��m����Y��p@p�qR��krh�McSJ��t�\�B���҉�)�Uµv��m��5�]�n����j�K�eJ^�+��n%t	f������U��Z¯X�����jsFL�|
_I��ϲ$�Q���0��DMJ���6�pK�e1�`KZ11�[G�I\ 3 �v��x��y��� 	Zy�����.s�0a��*�&�%�]U��Q(d���e�&��X́�R��ћ(J�K�Ӛ����	pͽ���p��ub����$���(�{À��r��ܯ���0W�t<�;�t�i�S�	x���rݬ6�P��#��ms�J$�*~��ωG6�J���x1R(�yb�J�BW���JiP�>��0�w��f���]E3g~�H�=_;��0*~���}��)�1H�)�9������am��Ee�q\d�G:��C��͔�97���
��ۿ=�k:k�3#tԦ�ffogE}s��w�8x��
�)N�۵�Q�ͽ���:���<��+�(H��Jp�LȦ^�6��ePT�y���F&�
1v������q�u6ե���0{�T��T��H�`�l�~v����g���tK���gvTC���
LͿ��%���a����)R	�6��$\����q`����D��_3o�U�lNʾ��p���eǁ��������B�郧�.�P��Q}⎑���
���P�3� |��9��8W�����W.}gwi2E~>���;��wh�(XĈ-�OL�Pn�3_�}�N��W�^�d�Y%0>�G���ɮ(��t�k��p�=�4O��{��VY�s��?A�D	I�IQg���L�9*%�������O97��7��{�߮0�s��8�(s,�ɫ���/���g:Vn0�^W�q&x��g�xԒn=����'	�7��jTD�	L�UU�pD��=����~%bHP��{)i'5؜�1�],J�W�1�#�ׅ??��B\��ښ�0i��2��L�[��F�cȕ�7Pj9nj�Mt)fܛ(���.J��9��B��l���f:	��
Eb�s�J�RĔ��!�o$��(��6~	R�b�GS�7w��,����ੱ����S dîҙ�,�T�ZL��s��;Xl$��6��Ͷ�>18�����;�O��7�M���s>/�/��"1���/�4�oywG-���{b�h�����`3$摲(p�n ��N��*1w��eࣹ�ds5�%E���7�;���ff��{O�����ǣ�wj0�aQ/���X�R��%2�óe��Ħ�=v��n� M�z��.����Z{��u�>D�?p"��;1��	���t�2mc�&�T&(���q�.�>�3�����Y��w�Q�O��)�:s�/�o�}��я�D2�%7P��)��Y@z��_f�p��"���խ,JŻz�r.������:��(�f���a��.Bfj^Z�cHAi��m�1z�%�VUXi�ڡ5�J{�U!R�<��[����������k��dY}�94����W����q����IϦ0�s�����E1�*�T�N��w��;,�/y��{���z>]��$��v�½�I�t�ie� �5q�;��8ХH"DD�����4\��W2�py��
6#��O�E���_�o�P�d�����@��I�JN�rZ��f���кGF�~/ŝ}Y5���| ]���Gǰ3�g�;l��f�Ϸ���ő�=�:1jxgO�>���k:��8��l�yYo/V�*�ݻ�H�c?nz�3/�瓎��t��#Ƿ��ۅM`E�B`r��c���˹�sи���Y���G*����:�Ȧ@��Y�w�PA�AR�HYp��DEǡ�d�2@_����s5ޔ3N��M�'J٘������"3~]��)����ԠC�K�7a2㬚0u�t�5��Bk�]n%c�H7� �I�*QR�+
,��?}��ч��\D�4�Ք��w���M���⏴��}���-ct�[�+	��Rv�����P��:/�9��O�]��ݿ9�G�p��qߏ9{
%EI�٣8��A()D�(�"�4~.�|�(�6B&v�V�/;��W��f���eqï�ɯ
5�d����Cm�S	��\Xe��}�*�_Nʞr,��+]�jb_˦��;l��
a*�g���x���&�\�y$#
W�J>�'{��#Mw� ����$�r��}�s
Ήz���da����{�+3Q]ӡ1;w�tL�kO���������U+=4=-�l�2��S}����f9ES�ٱ��h��1fC3n��Kݤ�����1`�'�lA�M0kG,یU�Uv�����+�
V���H���m���F6��.��j�(���̬r�h�3DIb#a�v��wgGo��mn/�k�;M8Qw�],eA*�ׅ�J��ˮBf�F��h�ki�\�5[sjJ�ڐ��sV�2����LbRC���5jˡ���m��J�uv˥����P.�h�G À��'uL�g���M�k=�X����rT΢�s��3�>��Ϋ�en��Hd~��D�`��3�|i,7�����9�v�T\�4���w�(�,��UbJ�Skiki�Lmcm�`8�������WEծb����/:�G�v[��fp����o�pA���=M&�����(U��Д�����O8�;.ky3*S�2�TL�4�):c��<g�������N�Q����k� ��7*�o�Eµ>��X�\��*ER��\aEgLLJ�/>�Un at�"�| 	Xt{]��%&"���XQ�#��<��L��2��'��*Q?��w����;X.,��ʏ>M[�����D��N{�xY��՛���	%T�C�w��gM��A��d� 
l���;"�	z�ZQ�,�k��dGx\I~�a����6����,t(.& ���D�U�Qam��9��[�B܂l���(����y����_J/_��U:�^J�v-8=�ai3¤n��c�*PT�CuUk<B2�߶"=����6o!De��>�գ���"Ϥ�5�(�G�>� ;�
�;�#1�Udd����PC L�܃�k2R�����^ �&2��8����8����a6D� ��/�;���-�Z����(E�ζ� �h�T�z�ڏ.׭b9^�ﰲ)D���X>���⸋��M�|�f����2�8V��S2�(����F���p��|k��Y�R�E9��H��?o�^�w�cK��/��H�O��c⟙"��������J�O�{of�)�$߷��
<p^���vT�<5DU.�c�$X_G�R��b�^BJ�d�F��ȣ�<��4Y�G��1;�V��"�p{��~<Q��q��K5$�~�.v�*eRb�GI�.��:��cY�m�mV�bX����g�����Sf�V,���C4��*��_�D׳*���_�|����>�}�=�W&���+F|"��x�<%��͇��~S�lB�����o]ɧF���9qӟ?���_��:�r)*=x�`��Kr�UT댑Ǝ?��XD8F�;�b̟�﻾��	M})��*r��b�U�Siit��*�r�\�E#��t���8���C]8�q�&k�
e�g�G�*����(��{>��2L[߯M�cpj�q9ד�����/����G����;��=#$6c�ENDS��ݛ**�-֛��`| ��[6|ȳ
���� �ؽ>D���@���M57�$}�,I<�d��S��iD3��40�<V�d)^>�f�ZT�ET��h-R�x�H�JfQ���n -�ʣ�q�`�л"����K6�m|2N�̾�0�ⅰ�sNH�삙B&��N���4\1,�7;il�X���uȖ��T^� ��e��I|�%4�D!�ҙG8�][��(�{8���YA��%��yn����4~�0BD)*L$i�4g]r���y����2�dIe�sw�O��]�e�qa�)}��pM��͊jB�I+(���
�ƌ�iu*Je����]�k����k]g*���|2�q�ʥ$�TL�3W8{aG��A0�[��2|.�]s�fH�g��:xz+7�y&Wޯ��\7+�X/��7�2s�wDÉȒg�bRt��v5�I���oY�$U�du]l�@��]~3�۴�FdmtV$��[��d�b��������1y3�uyV�]3�}8�U��q凍��l�>nt�F��VM+���=ݦ��&��W/`@���w%/deT��I8ycɢx��I�s�$J�m�SB!�T��â����n�GO
j�(�X����ދ��p[;�%��(U�f+]-	p|�4r���))BnP��m[@Ƅ%a�E�8��Keljf����>��|�mh�S&�"��(φi<~��3Q����5���싚xz@%G���іϼ͔�D
?"Rf�2a%o��#����}�
Z@tx�,�o�~$�gW9Zd�/"%����{���8c��5aM��I3Sti��4����Ø��fW&��������ދ�l�D���$�D��q�D*T���i�gˇ���� ���qF._بa�هن�ƍ8C� � �\�)8}G&BeS��)˚W�/z}����t�=�Wb߹�r:Q�[���}��Hwu;D�l� J��R���Q��5T�Q5P�O�v}���{wj��ά��Z@�
�c.6zP����a��ő��_f ;�85�舃.Bf��9�P��X&����1t5�p�GT��@�f�������4�J����`����
��ݰ[����6�tJ�fD6��bŊT-ad*���k�M��5�CWT݊�T�"KH����2]��Ɓ���=�XB1�p��]�B��cun�e�M��3�ne�.�qJ�WM5��ʕ��iH�&�x��߸��?��z�N���_�se^�ٞ�����7x(*ͳw(8���Y�)B;S.W4cX�5�@Ӹ��3���c��}�=��??=��&N�bD%v�b�X@tr�e�Kr�$�SK-e�ު�-���io���{�L�
MR�(� �Eg>ɰ͜ �Zh�c��/��K����oDq���r쎛J��Z^�p�9���%����m^�a��)�o�t��C��Xsbk� |ؑ��:�i�&�N�t�HE�gd�H�@qe�t�9q��Q��߭Q�4�i�n=t%|g19���b&��3~$Y��z��]6����h���}�A�'D3��u��+�<jWK��K�������䔨uR檦j�a�Q�p��TY�OUO�؅Q)��b��s7]�$^>��M���,����'����$/�Z�&M��ZW�٭�-�疄n�.֥���
#��o�<����Y���R���`�(2�f2��L��>������\��VaFms���4-���?���± �M��!�Fg?y=?xz+:��+�[T[�wM��V:�n�*s�#�u��(�A
�۹�BX#TV��2Չ��ͼ�*�l�#0��F��eYg��Z}44���%=���'�Ռ6��8g7U{�#�C�l,%��cHO�`�L�Y�T��&T�P�
Q �	ۧ_Y���n��l�w�6�̟C�ZM|=�>����D7+�)$uSJ�u�o�W�J:X���Yҋԗ$Q���r�_N�̽ɼ"E�p�˙D��i�jT�uSiQ݄�$�h�{y��,�tK/�5�;4�"6��25�z�"a���_p���:��R��R�&�0g��
�9��b�3W�¨e\�qD3�z��I`颳~���8}��2c�$d�����,Yf˶�ܼì�L���CT���P���Sz9��P�)T���uE௏���]�Z^,�W2�'�2�����>����+���� ����O~��KmJ����;�E�|z��>�F�I�g|�9���K�N����Y���S=�x��K��&dmm"��J�����E�Y����q��g����Y�}��0o�� ��'M���7��3��pJ��N@���f����Յ�z����}�@9R��]��0�sg2p�{�=(���A��3Z�a�~얱E{0U���"#4����=,����"��!���W�	�t��s�Q���ڼfl�+��5N�b��*�L��^�<�g���:�E{�z�S��Tƨ����"�h�x�r{{!S�c�����b��ק��.jc/`��B�FZJ��v��k)�'�^֣��s5TJ5U;.�ׯS�l����7PA�յ��:v2��D$�8�6C6'�U��À������bn�E���i��O��B�xFU*ȧ-����l��%�ۭ]�;ӱ�yNs"�կU��p�
���zj������y�RG*;�w˴a&�.���v��U�VU;�S
��m��*sH�$��v�]br\Vc�"n�m��эe����j����c��I묫�RR�}� �wp��ʜ�[��aDS�u�n�⡪Mˇo�UdH�n�?��ݗod>�]��2f�<�+o�J�o�Y�2����`���Y������B�n�<(�g��<�A�}>���#�6�-���z'�Eƅ��s1Z[鳎qm^Lr�m;<�&&�����]��$�>�\$`�~�ם����w ~볷��N`ŦsWvn���V��L��|Eo��n�ob��:7�5[�w\51�����Yئ�b�ofNr���"En�3��p�r/��̋}�茖W�d̼1���R�2(��{�q�/P�m\6��Y�}��#����	��PX>1N�v����m�dy;�x�w��a�y�������=�n����Y�P"֙\<i,���&���9��=��#�!����g�Hom�@���cf���=U³^�y��\ts�c'�V:r֋~����p���4e���h�5ՙD���K���3v8��r�n���Ntj��ڙ���N7�wt�<,�R�����}�ԩw��~�>�sN}��Ǒڳ���d&zz���'������śAo�eg4��5��S��;����|3N�'�TKw[��3�#lJ�_"�lG.�����<i��@�����׳��T��8P}�u ��銣1d��4��$����07v�sE1�������m��y��JIw��������Jt*vA60�k��6��U��M��LN:��+�O�cx��L���r��Z�����WGP���sU5�7s1���C�����8Di�q����a�D�ɱ|��>�!r��d��{�oS��ℍ�VX�ő�l���;��|5�n��`D	�ջ���=�^��8�a:��E ���T�Wywnj�KmhY�1�M1�QB;}x&9Q�C=�3�`�ˡ>��j9!��/���py��P��A��ݕ-�xfY�T����!�w����S�<�_�����s��.��*:����8p�霠}��ڐo%S|�)�R3�N%���Q��5��2V@������qj��X���K;|��L�}��>txV�}l(PM=��D$f�����.��YϦ`�?$M8 �2�iQ�$'�ι� �|�p`�6�4���p�$u�
�l��uWR2�j"�3��w�ei�t\3���ң����J)���:I�njmx���
P(Ϳ�ߎs�s7��Q-��U���ꄜ��NgӤz�@E���2`�KxQlO
3~��O3�B�?�!py�M���e���k��?6�v��ϭ�p�j���ّ̷��0�Ơ�m��+0K[q�,a�s5�8tv���C�+���o��m���]no�G��w��
(��w+>��|<+#'9��݈V���>3�lю���p��ڝ�SNisN�gJ>�g&�g���,�q&�o�s�������/�><U�^�}7�؅Q����5h��&GU2�Z��#	v3�s��p���{*�Bx�Ý���3
��	W��`�:l�ES3xQҶ!r'��'ۯ�^8=��w�QӇ����Fx�Q�;�{ʟ�h���EM��S'�ΦyNN��l}DtY�iP����Gq��3�2�H���q"��;����p�>{~�.���},ϊ9�+��'�+lJ�`�'4ώ�8�����Y�e+\�GM(({��(�Dk�֨ل��[H�ܧ	��[�Y11E�:��{�t��34�f�,^o���Δz�B"`6����tK79n�I��g	��+�_�g�_�O_>��䌧�q�Ѯ�0�6I�cS�<�KB9#HE��� �;�0���CKa����4�R���0VN�_tY���oT'�]
��l���}���0�U+M������~M���3�J���FotS 3f��\D�i���}q�^��U-�g�j>3S�T��˪e�Ĩ�of��N����;I�1'͛}_|�K(���P�����]���̺�j����2=�}�����y�����?F��YGa/2)� | ��=y�W���.�X�J�EuSiI�t��;�-aGQ`N~qEl5�]5�ϙ�#��QE��1�y��<9������*���{�
JmP�n�{Oa��]6��rs(���U��W�M\�W��t�ɟ�=U<g&Ŗ�/��<[R�e������;�9I��ãGk���h!W������э�h�O�|
y��CF�M��m�&w\��+�^�]�U:ͦ���J��k6V�V�X�`�&��nH�R�JvM�e���l���ιؗ���"c�V�!�UA�������M�6׶�^��0�, hT2PJ��ejdRXM��h���.[H��DԄ��� �|E���Or�_�j�9Ӵ��1&�t2��TLm����Dk�ض����J��2�"�����'�[f	�р��0-+���ĸM\WWL�kth��`��\2���d1���j��������Q�א��;p�!���Ȅ0HJE��ݽv������q5Ljd��e�Ӿ�:_v�;W�OaD�` ��|�����/�C����'K}]�~7aGҀ%�/���T���4���Q_dq�s@I�f}B3�$BD 2�����������$�	���PJ���eEV@���/�7m-�O�����%M��M�-��	Ǆ G^�p��y�<�L|�Q�&B*%*j�Hݕ��t\�I4��7�|2�����x.,uܨ�:T�t�b2�i��Ԣ]1�e9�0V��lJ�iJ(���Ŷ0[1f������H����pԖ7*{�������W��<|z��'���ǖ_�+��)�0I��Vt\9u�Aɔ�ʤSr��W8B�ó���q-Ir��Y�]̼�r؍0s���i�Bi
��q3:/ݙR����=�܎��^��ZME�ң72�r�u�+���t(��'Cߍ�0p�$�12
�/�	R5�؎"O��6j�|�m�ݪ�}Q>� ~ �.��v>@,0�>��q�,�g���4���t6uL �����y`�c@BfR�E)� ��:M�! 7�n�p�P�) ���y�_p����φn W��(��Rx�2�G�Kb%X�/
y���R?n�n|��{�RD�/!&�A.��c��кB�n�%I��J���w�r� 3[�%*�	^�q�
O"͛ݸ��;Ʋ��;�nZT=P��ǭ��������*`��h��rִ-�0Z�
J��Ku�|�A�~?2�C����H����Ň�5�L�G}]ʵ�<vP�s9n�آ"a�c��g7꾙ng���F��haT۪��Ƹx�*s֗�D4�D�Ĭ�?����X�	�nM�"���G3;V��D9 ��g��K�4�9���O%Y�C���l�9o�>��s���ۨ���>�QYr��2�&ԯ��v֥+��%�s��suO�X������\��o&��+2��S� �>`���qS�J�*{����g29�z)�[�HA��G�X#��+ށ���q�}�Z��7F�!�s̋���Jja���;;o�^��{Yxq��Oh֞8`�CN���h�쎓0-Q�JIR�S(g��D�O��^Bd"���*b:U��}͛U�ç5D8R%Bdn�[7��.�m��1���j��^(���&�\:|sb� +�nZ]��_Wp/ŖG�~ʿ�|�aA�Ù��gʺ� �������X;:�Z�����%Hi��w^��M��CL��u���S��0������4�9.ک���7FV�ҽ�Å�砜��Ӥ'U$�\a'��,.����aD� �@AN�vT.0�3@���@IQ��t�{{�};������nLW	4K�>x\;;ͫ��G���Yɼ6"�!@f?��x�������|(��}4�ħ,�(�uU7�ƽ݅�/ĭ{����4f~o�a�,�`lz�0�W0k�G��oojP]�h+��7����0��`���;�?aS�4g�MÅ��3�l?M<|�{��r���x�����V����%�S�[��ȣ.��x#*r�g�#�9�J�^��灤�3jǍu��t�QĤH��ս{��C����b4{�y���ܧ�W��Ɓ0����õ}�_�],s查����h�	�W�������IㆤDp��߮o�%�a�]qZQr�n(
8�H�������,2�v�X�L�R�,I�:�Ic��i�nT�͓�������[F��PAʲ�ՙ�v�|%�u�}'��\;9��_'�Ku��u݈��!Z��5d���h���ۂ/���R���*RF��>[��_c�H�� %båo׵i3ŏ{��x�0K���*h /�b��6��x"I��_P��ax):X���WǇ�9:��\4BBǟ>��U�0J�;^B�F�9�ɠe�I�S�IN�آ9xC B���v���m-�VM�Z5� ��b�>�����
�3�k�.28QS�#�H�	y �eW�2qŕ3��ߎ	V�IĀ���wg���|Fn��`A�R��_"��>��ꏟib�z&���YYAXm�QQїUϬB`6����fwr6�Oaك9��>��~��8c�ǋ<�Y������[����S���o�z�G"��t�cv,t�՘n�6�Z:e7!����e�msq+�H��uL��T��uQۋ�7���@�T�֨Z��::Ẽ�έg즬����XfE�`�6 ��Y�+c.���e{[6�I2׮�h��f�3.�k�6�I�ɊƚڴK+L���Χf��mZ].�	tX$%�%�U00fL2��p�����|�<��V	��<�ri�ZDC��ܘ��ڡ��숖@��
&0�Ɍ8=Ɂ�F*} �?/j����8�+�%íŵ@�&��HZD5sB@�H�i�Һ $�sp@�;f�M�u%�29��H����U��=/��^;��/K�o3-?�I5ig�u���zJ�K���r6��)���˗~(^,�e��6!�@Z.�M�,�r�&�I�p���W�(tP�F&�V����J�)W�#�����N�#'^E7b�$Р �����Ʊ���7�I��%�șni��4�x��bO�	>���:}g&��i�c��o���+���T� �	߷�Z0[�g�Yi���9R&�o-*��w�W���w���� @�����S����^,�g���8t��]ԣ�|v�3)�e�S�r�c��,c^X� �4�dÕmк,&����@�I}�L�ff�f{�'�=5��'Kvp��t�+���#�1���~��W��?�R���&�PQ3T��(�������Kl�[R���������MT���mu���T��b������nF�d���y���*ɾT�~�>E�������X9�*ï�\��^\�L�X�R�.]��ڠĉ�#lW�� x\!v��wK����õ�E~��Z��.�7����A ^M�܄t���Z� q�3�ƴ��P�������άڦ�UK���i�����P�Ǿ�T�a�B����Q}�2��3I.���J�,�����g����B��%U���/�M�� ">f�W8$c�s���W�Y�YQ�ĝ/a'������/������r75R��'@���ϛ�s*�J'��؈vF�o�����n�+�S�����]����bݾ=����*D&��a54��t�V�c�b�K5# �٘K6k�v�>� 7��A��s2�nh��O]f�1x��tj$�gk\��=��A�8Y����L�(P�x	�Q_``��x�i��p�r����'	/������	aF���t�=I�4��O���x�6��T��ҪrԺ�/ŉp�^�^\��L��W����G�,�󣊮�}s}���D�ȝ��Le��!
� @��guB����7[�C	�/_co!Yl���==1皞��&�.�!äV�s�#�x��&�\=
�Jː�]��;�����F	�ZA�)cWfğj�N�cJs+7��O�Sθ��Ό����x��G�ӜS&��@d$�Y =�x	�D�H�}Y5�]��-��\>o�'>���%㏶:!���ٮ�ŧ}�x�ٚr�M�4���%'�7�x�x��8��@�߹e��.���~<x��9ʾ�Μ=;gƶd�jٵqmIAɅ���dp[�i5��2�l�i����'�޷Y��9ϓ��g_���~,K���2o�:�/,���R�G���o�,𗴜q�5DL�fd���/L�"��O�3x	� q�����r�F�ن��^Yx�	�t�I؈i.K���=B͕-����7S7��E�����"��O��2�b,z�N�B���/)����~G�x��s�Թ)MMUW�Y��DJ��;M �Q=�kM��w��d7��ں�2k>�����W6�����ϣ��L뀎0�����a�����C�q�I9�����_��f|s��C���O�$��O��O�H{�>+/b��Ng�lсWU^_���pӳ�q�޲8U<sː*	��a��˝���|<c%�^�<�B�`L%�1*(3%�D�)�5�� �xH,�3j�C���s���=�-Ϲ�����/^�W��7ʢe%�S2Ы�X�R"�2��n5�f���֣^,���`}w��JQH��(���x~�zO��ӈ_�7�$e񓹘sT,pGXY$|{w�;�_�╣�.!�"�Kc��~���Yʵ��TDȡpe�YC��*zx�B;�n�٧ a֯�7��{��X$��GG7�v�p�.����7=��b�,�0�L��{�C4d���X|8�CS��q�gM�1�َ�3T�J�UU5�t��
^�Z�9�/K�z�κH�+{�Ң���E� H!\7w|��rxKp�/�8*A�L���t\g1_��QuB����E&V:�(�<i�^�I��r��]�T<;���J��N�tѣ��-���3l	��{���d�/<�kH�!�k�K��G�K���Gˬ�F��Y��G��,��y�s�\��;蘣=X5��cLxnq�餒�+N���Q����D+���*�j�X��btC]i�b���t곕3�s�����Ǌ���ɚ<��ը��v�:��aB����,J��wYJ��n��OJ��pt��bRI��zd���zw?��5��L]M���������.��Q��7���X�J4�.�P�|��{���.&vPYW-�:�淶0C�AF����ױӚ.����=}ʢ�"z+C�F��;���uGF)Y{���'bΊ��yƼ
O~�ӈ�yC��r"�RK°u�$�I��zEr��f��ϊ&{��H�{< �>>h�7r���Q&Nƺ���/I�\�g*������+7i΃�4˻A�T5��D'Hf��k�v���Q�q7b�og�*�]�Qh���qپ�N٩�r���[����k�S�s��Ù3����s ��*�.���3�����5nCH\b��B�M�Jc�k4e����G;��w{u��mfN����.�6��Cwc:�Ȼ=�����W|��u��W�zq�Էb�'���R�~uR�2��尿+�v��,��4dN��^�g�{x���F|�rN��ϳn�,� |(���/Q��z�_�+'n���c]�����KSy9�Nr��=B�Q=�81���MZv�SYyq�"'D��g�:��I�c�z�2������W�O�^�����)`q7�1��T,÷������}�]UT��Yڛ��Dm݃�!P}r6ظVO�o�rfF�рΨ�b���0*Z�ye��X �	�u]c�e�:�u	��Yn՘��2��Tg�d-+��G$߀ �E��VX�L�N���`���
.�*�3z�����eJ�c�),U�0��v��z��]wb���n0���]6�.,w ���i���WQ��]f�B��<e���2˪1����r;�!����b�)u�l��xλ�%Ꭳ����4�,`I�LkK��d���S�r�,j�f��5�h˫�lul(�ivt�t��s����,�Z����Ĩ���Mlf
���Q��5��+t���䕎��вZ���03Aj6l;� j]����u�U�.56�,B%���iɠ�%��0e���é�Ļ\�6�f�L�̤bh��,�b��&��vKƉئ���\!��du���+��#�ZR5̪[��h�q����Mc�Z�f�����5ٌ)7]qi�<��4M�I�MDm���Q�Wj�ͻ(�G��[7:�h�,��(݃TFK��8HK�f�퐲�/Af�SBk��]6�[F�	4:1p:�H�eJ5+YQ-����6��Z�H���v�ƚD(�"D�b�W[��H�J:gm���0YWqvb��be7U��ĵ8��6�x,m�z�5��Ǘ(kf�*d%�Xv�+�E�q6���mBnL�5��9m�R]I�BqHV:\a4\���
�[�mԴ�#s���ue��7XLgB`���2
7�]`n� A��pkV��-oW9�F2��2�3KcT4�LҶ�莘iI])m����`�@6^r�]M��4ʊ��P��GZ�	@�u�����Ԕ���{6%1� �jՆ�X!�B�	4�J�k�]�)Cb��U31�
�sd��ZT�kZs��ӡF�Ŷ�y����][�0&r�EYu�.�kR��m�H���4�M���PZ�Иq��l�V
�($у�P^FmZvCZ5��ch�m-T#�u��Z1Ym,`W�)^�DD،�m���mA�C��Jh�a��q��X�۬t��D����������g҇f&!IE�Zs�ph�2�1����S`���gi��̜��\��
��S0(D�ަ�v�;��=�G+>�ʟ�o𷇁�����U����D��q;�Cy�1�X�S��n�j`fe�ڜ�ݡz�^�>��k&��JX�R���gk�/c�j.�1�S�q�5fhj@���J%w���m=*@��_K{.pA7|�mlA��`���v�cRb��u55���bD��N8{�3;�ERqC�c$�\s�w2�yQ7��pWtq�̊������p�(�Y"�[Ǥ]H4cu�PC����cˣxoM7s��r���41��r��M�����N���i���Zd(5V�����`�0���t.˳($�&e�(�̨n��!GŦ�9�z�z*"�U���F����@�u5<�
��oGU�w�u�wT��+"T�]a�u�Y%����@������[l.���HL�4k�6�q���sJ�-[�F#D�Pcd<���v";=9IR���ޞNi�`���v�"�Z�����hＳvx�S%>����T38M!u��;qz[���w�쌱���3z������W����H���>X�Sw�d���r5���0:�J����ý;��l�[U\x����������ڎ���n��noRj�����g�����S�0/��B������2�4j�Hɰ�3���9�7��}-l�aSQ�q^VEh�ʱO}�?uЩ����f�!I�&�6�F�H�S9��r\�k䗉b�ܻ)�4X��n�F."�Z6�YC�qJ��4� =f8�0K4 ]H"����Ӎ0�b�(U�`s�Z��oս[�6��f�Ю4l��f*���R���Z�5�7��dF�e�� �$ub�%�kM�̀�W�[W��3M0#us5�M�a��#{���\��d˧Q��xGd8�`�[nzN��Z�o�����36���W"�؎`R�;�/q�ǒ�/3�7��j�@���)Xi`,I��k¶)`���U����ܕ��i�6`���~Èq����B
��xI��)ϸ螓�3���3�$�p�ו�8R�O
M��|���ge�$�"ee(IEqx�=���O�T*��B�âݯ�7҄�N�:IU�}�h�� /��?D�ʜ�L��
��ZY�)��M�����}�b���4Ȁ��6���@�6{��g��f���Q<%$�
%�+��=3�L����ӂÅw׮ң����kS�?V�TZAG��-2Yy�0I�9艑2��J��.�ܼw�5G��ż��q�/�x�[����͉Y��Mt���6+�Q��v��<Q��bV�5؛�]2����iRV$]`[2��!GƳչ�6
����=�_M4Y�p�M3g6�}{���z�-ɔ������1�0�{y�mL�IL��(��d"͑�݆�> ���#�����\VD�i�w�O��grd'2R�uD�0UUe)p�:�
�h���Reh�%��}r04�܊6E�0��3 �I/��ʭ
BMd[�հh��l҈^7C^;�}oSϏw�Y��=�ILh:���^q_�
G=!��}�wӂÆ_��������Q��@��+{ �|���T�$�T�u߄�|<����G0��$�����Qf�nu��D�vϳ��'�b�f�{� ��7yE�F{k~�XI�.ײ����Ӛ�6��g������NQ��J�L����
N�
}˘��:���� ���j�,���37�7ӂÈ������\�P�3tsM�"\���L�VZ��ciJM��.`a�[t��;{KU��~wO��fP4�����gP��g�c�B�:��L������RH�B��F���r7����W�h�2e0�UT�t�+=��̈́���Zy���K�q��udP�J>]4��xH��3���׭�LҠi��w�ZQ���'���2h��=���q�ʊ}�ww6Vn��eY�k�������h%���Y(ߛY��|`Q��j��T�����B1u(����*;�ə{�۹v$I�\>�k�r�x9�!�������~ݛ��Ɖ��xݿ���|:��~؊��R-��!:��`^o��WЏ��O�Ѣ����{f�]�͐�	Z���c���H�T�*;�CQD �������	�ea��5MS>E�G ��'w~w��ţ�b|�:������s5q��E�/׊�Q}I�^�ォ��qd�$���k	<%{
/������4p�X�U��miqK���k,hK��Y4��26�y~�;��v��֏2�o���\1�}���	�ԫ�����n.��sa)K���M>��}w�;�>,�ߤsәةS%MT���^g�=��=��qC�E�#7p��A�,����O1(R� �":a�Ub`�UB��*joEgK;�w�Q~ci�{�YO٪&) �x���+J;ewfғ���ɜ�XR��d�M�T> <�oʍq����Ƞ��{��it1��=�.3D��]s�ڻqz��J-�����_��[��Ხ�r�P��q�O����.���r�Cf+���=!��(I8-�p���P���Pj��d=�ZŃ���1o��2|�_�[/Dzf?�_34�ov�����P�dLq���Fl��t�$@���Ҷ�]��#��A7���)J�� #�O�������E�3�W�W�C��v��0J{>U⏅�R�ߒ}��v}F�!���K�XL��lڥ	ij��BnP��%Efŭcl�;�"����5eBJ���ﾹ�|�4�v���Q�pY9̫�����/	�Q��U��<|/��%����I&���B,���UsӪ"�E�Z[��M�'�����ך^,̫ɼ�*bRDl�}���Jx�a�`�UÞ���Nf3|��g�|;�� ��(��<s*������{�qe0�#0��4��&jfY4^)�ԑ !t��y��XY����~8M���
�̈́�D1U��xH�����Ԇ�M�T�����&Ң��s�%1 G��j��bδ���ߑ<}��gK�,�ϔ-Q�?9��'~�o�Xw�u����Tγ��dMt���#�N�,�N�n�G�E8�"#�������x�R�Ur��lU��#b�όig�~{�6V�!�����2؋.tֺt+W�-�b[\�n)���hŌt��GA�����X���+��é�F�V]��Z��fUF��hDrL��R�K��cUj빘�k/Q ��M)��.���Z�D%�W٬u�6\j.�ݦ�baJ���"�-B��,%an���&�m���bD��6�(�.��$��_���y��z��"����
�Pȍd�YRv�]:h��!�t�+� 4���~S.�->-܍�+>@��rq(�'Q���nJ�Q�[+�f��M]���A3�],��F���$��4���J�⢮����?�X�vt�Wu�+�v%���u�jPG@�-:,>+9z�H����+^��Kizd�T�:@�.6����A>$4F��yT��N��⻠aw�]u=_ޜ|���~1��Ԕ}1^�����Q�+K���ob�]� �xp��y�f�`|p���K��8z����r�h����x�J� Dpy�;7:�0�Z���(��*Sb��>;�ޑ�#�J���w��å��X�t�0nh����}��}��XQ��L��Ӫ���'��ɾc�FVro¤t��R�j�"֠p4��in-즳%�-�a��4-��8��j����o���;ٟ/���]6ɲ��K����@쯰�"Hqk+M��-;�_1/�P���g�ɵ���^��KA�T$�T��ӆH���3��T'>�a�+����O�h��eP���-Y��v�}�<o�.����d�+�>�IpB;/���5�5&w5�,����z�-�;o[�t�G��}J�<�U�?�4p�Mכ���F3^jˁ_9jǮu�8E�ʽX�M)�w�vR���HU0q*�ȓ��Tm9��l���ؿ��\A޸)�6E3"l*����ޢE���{y7t���gU��I4�@�U�N����ټʿ�_-߯~~݊����wϳ�����OB���3K^���+3��](]��B��o��w
E��;�J�MK�jH$uO�
0�+�X�t��_s�P�I�� _}�o`:W�����;�<<��l(W��k�#i��P'5���"U�Cj��^�*iMx�2�0�`�[��i�e�ha,d��ҷ�b\*����$X|VVd��Q��s��W݈N.\ Q��D������ܳ�T�*�U[�#�����sb�a����u�vF����E6���yWN{a)K$3$��vCQ1"�
R�(�6[��V������������-�O��������3��]�f�����'3�3Xy�n��g�Fl��[z(�G�)K�w*����E"���{vG�����eƭUmP�"Z�듸�׈X���z��W��G�~���xb�0~C�i�Zr&2>��kfPw�/����#�mv�,����s\El�6y
�&"҅0�2���}�E��D��_&�l��~���0� |W�y7
���!
HK��Ǻ�h���Z��C�3N����p�W2o	a�saE(��9�[7�����ٶ�	'��q�^q^%cz�7q�9�r栛m,b�0%�vTM�ԕ�]�ڧZ�&�5���E��v!;�q6R5.fi^,,u���gK338�aG���\}�V�C��	J����w龉aD�Z1�P�̢I����,�����P�H��yW���.ww�8/�s�eZZ��! q��U�l�9��R�eT�����"�R�E?qѷ�L�~�� ?��n�o&VW��	<Oτ�9)��"fhs.�_
#��IB�Q���.c��9��,!�(�{W�Y�b��}�t>�ڍ������2��y�T�'�y�$Ib�{F��ewt۳&H��9` �@p$�r�X���S��y;��'��N���j�$w�l#v����S~G���aRs �S�&v���j8&��X5�p��3��6�d8짂Pƞ�ɥy(;��E����>?��a�$���[h'A�*	s5R_�"�M��w��e���Jb"���z�|Q�<"�|j�E�g_�5��,������+H=v���ǐ�	���,��&^Yb�Z��D�B��*�t�8 ��i�WJ��ܮ�e��@%�R���(�ב_BX%��6�o'��rxm6U%:e��>��0���3��̈́���@ ������#����Ql�F���Xg>��<,�$��軼�)`�*�C��/e��|?{{7�.����7����������q�(�F3�i�:��*dz��4�Q357��sT,�� I�i�����4a��(s�0d���2��ԓL��|g�ܛ�K8�v��4�t�K���Rt���eǱ�a��P�(A��گ��溼ҼY8W}�w�4t�B��R,;h}��!�r���;:ASQ��"�(od쥧�7Z䉉��ȼ�Y�Gt��c��|J����Rx�~;��fZ�nȒ�q��k�%�]7gHu�yjFlɀ"�]5ki�j�1�ؘ3�],k��P:ӡ+Ť�u�+65��əH-u��3��.0�&�G]u��b��H�ݗ]�h����j+�Hع5�c.Ѧ�]+�P"	�� K�C(Za�dj!�Q뺣��m-.y�Գu5G"RZݐ�e���)D2]�J�Lfd}�oz޺���!V(����+�b5,��������S�gx�����t�R�+B��	m:�o%�Q��n;|�Cj��z�S�ݵ�GV,Ԫ�%z�t&0�n�%0M6�1,Hj[L���I6�I��m�)X9Mȳ�=�2YQ:�f�
9ٜ�y�؅)2�/�(�:�(��}�M�TB"fQ1*P���q��ء��BIw�i�;F�Īߋ{�Z��~����<ԣ����ڴY�Kژ���a)�@�f��\E��gygW���l(��Iw8o��W�Ӏ�;�U҅��G�ϙ��f@n\ӻ"��D8J�_���XQ����z���g>w�/��
¡ HGݿM��òj/� ����kp���䆌���Ng6!4�wٽ�Â�Ƴ9�iQ����XQ���Ӱ���q.[:9C��t�Ma�t��j�M3q(�Z���Kp�aH-"P�'{�=z�_=Q.Dܶ��t��P�/����x%����9�|�,�yj~؄�.�"4�-gʱ;�e}܄LaL� ��S�,�]s^�WP��e��zl���Y�d���V��,����[=6 �.����"a=SX��x8����Vf�����\�NL���{M�j��j&w���y>��ꑾ��p�����>ڃ�d�\H^���{��,���ɨ���q��ӧW6����F=��	&$�aÝ���t��]��/�1�]�8���
��F/lF�'.YJ�A�;�K0�~{n0��_Vy_K9�� ���~ٽA-ac��fғ��ȥ�bX�Rs3STqp��
D'��5�����Yz@g6'뾊�$鏀�%����q�+�w>oXL�����B*i�(�Dbl�4F��z � z
��K(���o �ǈ�ys}(����b#۹(�F0����R�T���[13�jXb�R	pq����D7�?}8�򢞋4���޽��?n���Qҭ�^q��vt��/��W;DJI�
G�%���m_�qM��B0T�0P���)�Q���\�Z�5��+�){.��,��k�ʿ	?>�ϋX/�!\�%�ď��S�*�ITR�ƌ��6^�|�ę�x�w_�TO����s=��Ev��*�T�D,�A �MCB�"��Iަ���w����"=����\���6�o�=^K唾���!a����Ax�
�Fw�t��г��$��F3N�*
�c3*�
�",ho]���'���G4�ʢ�LOT*|R�Y�dۺa��wJ�����1�#%d;��D�T�>Nlj��Fm�F:8ܚw�0�>�l����`��5!���{h�87����\b���q�u�qS�f�rfBg(�0��n��QGu��F+|-)#{R���I�/�bΡӛyT�L�p���{sn,eo<
��t8V��,�l(=O���|yJ.[���\(�]g�τ�{���7�
=�o[u��ڼν�<4�m��߼���$^�w�Y�x�w>f]�����"���s�_�n�/'qɭ������1�/_���T�|W�.8���*��wU��ˣUUԪ��6�U��MT�m�>�IR��9X2Mv�MLJʾW�׎�0��-������=�%��'�C��>�����W��#�#�SW5[1��J�I{y��gc��j1s�gݓw�1��?~�G���\G>{���u�QGj1nv�)��ޅ�����'g�<��яO�]u��v�	V{.C=l��Gn{������Fm� ���	ƞ�f' ���_�:U�zx�����*��yM�z^K��y8�xaۚ�6�5p��&�<G��aq9�E(��J-CN�^�nd���p��Lr.����R܌3������=1�
��~ߩ iA�!�m3s`��l]�\P��(���Yڜ7"����E������"��-����?�wp-���!~EW�t��.-��Q�*&Z]�������$>�9�i�I-xo�w��e�;v8����];�w��1��ZYْ���U�ӗ�ޫv����ǖ��6�+%�c��6kz&\�q'{��]���A�$߳�@��[�W��\d���k2�m^f�/#kr̷w��6(�Vo�)3�:��9��w��\GU8}��c�3k���8�\:/������yA/w,�Y���^T�{�.�5�1��������w\UN����ew^��C�C7������f�/%�u�TTD�{&h_k���ꕪ����c��S^��j�xM8��j�r��#v�Cʧ��>驵\��1w���7����7.@ª"fw��V���y������Bo��.��x�dM�-�V-^�WE���m5�`d'�����&%�o��&Y�9�g�LS�cs�X����>ȗw�����ܷ����ػl7x0'#&}'%؁y�ĳ㢾����g��s�G�>9��ɽ�Ii��C5��1��ڙEӊ4m�Efκcv�}\��!�����4nM�MBu�ʻ-��U�[�[��mCc˛��������8���C�ly/��>�}��M�7��O^�D�-�yױR�i�\��8LJ��m�`�N�nr\}w�-�2OI�7|G�#~koE-����?z�f�`���g�g����;����������1�����>USU/t+93�B
���*���{��1��3Z2l��(+X�JC>�TݚY$�DذP���*��c�|O\q���6#M���48�ϸ�	��BjT��N��J�ГR�I)t�����,({��x*���_^[Vx���!&�.��gد��G�/rީ%(R�T���8�œMu���ܜ�@|I"������S(��Y��j���� ��O�|���RR�ll`��;fX��h1��n��h�֋,�tk��]4��z��Ş����>R�����6zn��vFp�:�W|(��+� }��¥�E�ȝ���UCNfiP��T��;����jP�> DY�O�f�꿄��=[yW�I���=Ix�����	�*T�xç7�Qi��< ��o'e����
���&��I)��,�Nwj�0��b�x��bqG��`�1�D�����Kآ�S�����ָx�&�-Y��q�W*�\d��<+rڂ�>�j��rT�:~njG��̐:�NH��6�X�l~r*�lR���:e~����dǛ�Gxj�r�>�}�����)Ѿ�v�����IW���f�(Ve&��Pn,93j�g�+f.+F�����3EM�����L>	��e�o������ V}�<��x�]4���N��ni�|P���^s&�t�JI�-��v��^k��w�	x�ӗ�x+�Ӈ/�i��}�-��5��KU`1:��Wg%!� ۝Yv�*km�a�mK�_N��:+��Lg)�9���4�N]��|�\0�����xH�Z32��+ڒ���9���<�Д����L#�N�e��5�T"1, �d��f�(}��go.0?�\��+��N!+]p�OܘB�vF�neә��Œ�N�q��(����V;;{	J��A6g�_�:2����_��Q9�V���:�3)˪�cVOoR���"K�'H�I���'=��"GO����x+TD��B����Җ�q����~d�IPB�))��Yd*�d��_��� �����g�g"W�sTYt���u�4F1I�=��?c��b��$bۗCm`�����	�*�,Gj�5J���'���s+6�VpjBV�Nf����i4�σ���N�`7K���S��&��u���4�;hv��Ʊ��j费&iΨڑkf��&n�*)-(�mX��4w\�F8*��7D�m̍Ict�/^َ��A4�Zt
:Դ.MK�b��yerK�V���m�#��@1e��b�	GF�f6�b�L��-��
�Q	p�Y��dM�u��Ҋ)
��\�[Kks�W��ѳ)$$�����#��:ɑ����w��ݸM�-X)^&�3��s#������9�]��!��~����=ĠmT.�������Xs2��Ж��
�t�lՍ�&�զb�]��wMz�5A�$D�$$��:��p�})�!�1�睤�Ҋ�g2y�؈��BTp%��6k>5�H�*�~"G�LL�$��$���ӗ�x_s��L���;Qg
0�.b)�G���d�l-����z���,�ี/A�R33Nғ�
��vx�l>#�O|�z���$ 藎Q����K��2(.�C%�T��3SM��Z/�ڒx�J</���Q'�^�Ҵ�l�m�Pt���O��()��x�i�i�F��9(T�C����6p�;=ة�O��@A>q u�T��C!I�@3&͐�6>�<�;O��_�y�JF��9*��)��Gk)�,6��:��F2�Ϲ�l��g��dJ*����M��t�s~��T�K{�6��	�O>��(� T^ő��WEtK� ��	S%��+:X��W��5P���W��9އ�����z�̬I�Ԭ���_��xR�~Z1�T��>�V߫?}�x��V�o6���o� �����q��F�U�������~��������L�bXy� ��a�c2����$�0)=6��tV.���� ��7��(3$
;�қ��}.y~-.�C�AnϏf��J��-#��f���F��ye����3���_��Q�BKfN�z*<Y�^���3�a���a)���
m�����Q
)	t�}��|�GL/�~�|�)8Y�ﲭx�~�P�Wn<ϝaG��v�Q0:H�J�S)#A��,��d��J��T�椔H��{�Y�j���xM��/��M|*N����K��i����R��I����Aͬm��a`����[���$	�oW�#κ-�o�}	��ɵ�Vx�;��WÅ������("��i�3W�z)=����R���S����K>rx�Wyx�O��pJ�I�"��2�_�T�����^\��D�mSʵ�jX$ؒ_Kv�s-��rR����E����|���2+��[y�#�u\}�:����2_+�<8�>��\���7k��B,��{V,���}���q��A��1�l�5�C��j��|��ǆ�W�'b6�v���W�Z��2<���҄��� T��؂CD���h� ��B+Jڥw�����I� �A��u�(�z���
D��K̩r�Jt媥Nf�Z�5EBKD�x����)ǭ�;^ٸϝ��y��I�3RJaB�{�vo)���05�e4S�C��x�*�9�藉<|N�'�D)���.`[I�����8G�E����(����lx�>RHa+����L]n�XH[Qjd������0yqe�&��wO��<|���9
j��؟GSn����Y[N)���s]���a��}2݌w���J<o�d�c�j��D�*sSxI�k���̈́�%���x�s�-&xᾭɵ���]b�؄�%h\�I�jN�h�rJ���������Q�r�����͕-��/�z=�GF�k���b\'ٹ7�N�:\מ)T¤���T��L]�vTG�Ӟ�굼}����Vd���n�M2/���[']���^���������w�' Y9��F"|����?cؗ}�;�E��4B������Ҋ/�>��φ��ѵ�� >�n
@я�J��}0��{<��/��Z����Ô�t�t�޶{{�ў��?�C.�8��>���˵Zd�=�jOL��[ST�MM\a'�//�"W�j��`%�sf�T,8=���)+�ŹY��������矯_��l���-�\�	�B�f��
�˃�l��n�+��~B�w:��)��H����g��/�ɦ@g":p�(�����G��{�@eq�R��3����L�=((��2�YC8]:�^Ǫ"T$ĸ`�?}��ig�R��^$��|v��M��B�	�R$��kZ1�fbW3����w�q&͐��n�!&����zk5ذ�{�b���4���K�b��lhuSk
>�DT%}M�oE�z~�U�aD7и�F�
�P�BV�N�������&'�fP���3FH�d,��S4C��������zEp~��k�|�*}��*~���y#cr���zNh��'/�y��)�ۜ��O+��*���՜5��O�A�g����~��\i���D�Q�
�n��"$�`�BfB[YT�%&ۊ���]t���\6�l��DR�f���
�.k��J��@�-��.ᱱ�:�a!(�x�c��ƛ�3$�XŎ�R���ae�Vі`r�uI���f4mH"A4�+ex+)��ds6ѭ1 ��3���ezۙ���S.Ɂ��P!��-W,��k����4�BP-[4Ys
SC
�]�Y�Hc}"�8�ӟ���[���n L��z^x�� �wx[J�k۳��q��r�{m�R�\o�Сc����o1�k����$���	i��cf�u��1F`l1�����eһl�:8?gt�;�C5��� [S��y���S�N�W^�ˌ(�ς��㻙ka*�BZ2�d׏���O���rRs4�"N�V׳w��	\G��B�P͝�c�u�@����'b�cFl)">%𰓛�8ԍ�SD�
i3 �D!�W
u�g__*fJ�Bj#�,*^l���2�r~�����tj��x�@):��N��' ݾvm`�K����W<*Ǉ7���6�F�������ó
�6�d%�ɡ�ߊ�}SYy�Rt�{��x@B�o�����N���p:��=ϲo�B�fl%�R��̩$NY�H����v]R˄�00,��"kq5Kf=t��5�B� :mT�2�oH����Ꮾ���ئh�n>}}_xy�ƈ㧾ynҳ�OW�
a�(R�Hi^��EOY]����/:�w=x�i��ed���&�4\{~x!G�+���}��H��uO�U���gzD�2;[q3W"��z2v�Y�X+�Tt1��D�J�o�׸!��s�_�ܺ�ut9��k8w���^�6M9ܪb.�HN��j��r)\�������ed:��V�@>�3]�&��g`Asݕ�I.LDE�p\�6�PMM:u3U7�H���O���	��������D J���뵧i�kkU��'�r���Ч	lsH%S�57�=��QI.	%�+�V����F��b��~W�Ĺ�RR$��BRz�{7����q*u�M!�J�M��,fb��`�㚔8Q$ O��P�.2u�ˎ��d(�o���[6�a�N�UB)N�m����P���5�.�v&���v�&�R�m����:@�?T�n6�E �i�����|��gƸ�έr�9�48�SnlU��	�	 +<.���ŭ��wq�`�49��ST�����9�~��H�0��5S4TaEN����8*���~�L�	g^O���S.�J�5PMQy�m�Ʒ�|wdY��3�,؈�9�*O���rij�?mAU���k[$�R*z���Sf����l���5��8:��g��֡���2	�E���>�F9����/��bA}9���s����&>��F7�TLD���2�l��Ƭ�<�)�[n�/eL�ء��)��6b~�>� HeET2 �:ɦI�GߐL�mT̪b�3U�
��؈��@�(A9�6�Fab˭ʾ�����U����(Q��y�+Je�fiK�'�j���-S�v��x�����OϢ�a&�D�?�z��_7/U}�Y%�9�K�:p\�̈́��xk,r�:N��)UR��@�Mtl-��&�6�F����h��~zN��e���LL�L0��h�g��b�q�Q�8q*K�ي͈MG��%�đ��X��+�O�k����S.uR�.jo�_uٔVro�jP�E�/�㯝gw�,����k��,��2��u��=�>��A��^0���L�iI⍟{]��̦�L��MJVBK������,����q��ȶ*����	�R�U>��z�^��#����V��4�'w>w���<��J��aG�{�����vsM<�5Kݚ�l?�`o���_/
2}��:D\
�2��(��/Sp�#���_[�5;f�+q�*g�0<�sG*��.�L�����K�`G8O9v!�t	3k�'P�� �zf�c:�!NḰYˊ�.�U�A�.��>���oh��*_D��$�rrI�I0ꪥs
(�\3�}�\����}�D(��}7�)ok$��Kf;�3��V>KI��lbh�����~�����v��Ln�ѣ��d���W�%IfBY�p��I?$����ϟ�r&�nQǿE�N��>-):z�Vg����,��v�!$҅��ïn�s�X|m�#���34�i;�2��M9�T{aCP��@"Αu��k�,���Q�u�j��ڒ���%�Κ�oa��ӗ2:t�!CM�N��!"�묚� .��H@�<afUo&�.���֬Ç�����|uN��TQSN�Iͅ	.O'���L�������Ae�|hqD�o�a.
ā({�[�(�n�	���QI���T�����=�U��şlBq(��ֽ�6h�u��� ���ɦl����hd��f'�V��<[5}�qkhJ��?-ō�}���K�u�"�w'�uy%��o(I��Ϋ�l`�a�z�Z��S=7`�޴]ůy1���ݷ�f�<��5��I$j8�oXw>@���fk������ �_�O1�C���bob�d���j1{'���5�j;K����&Io�?gw������M�w���x�O�Q5\�vv���2O\�:b�8h���I/�V��bgp�YOt{�����m��w�n��E�������/]�v���o�c4��;��Z�{c�݋�zB���_���3�ZR?<�ߑ�w��95^c���:�M^�;-�;)����.E+���tD�66��GGp�qם�ƙWlŲ�M�eTؽ��N�m����gs5�4��9��d~��l'�������ک��<�P.����n�T����!���j�2�8��*ܮ�,�[��]s}��r�Zg�G����yFy��m�Q��3׼���(,�Y�&%8��lXF�	�!LM��k!z����O�w 7W�ͳV�8{I��S�<*aE���=�ӝX�"DȨ�&ZY�Q
:.�}>h+�~x��G�4�u�~���
�=��(7˼����3_��{���u<6����O�
�g�}�d){#�1��!��J���!�?���L��W��}L6.�~.��s���@G� �l��Lpǜl�;%-r��4u�FY��L+8���p��i��\�ڌ4d�[��l��Uכ3�'d�B�j� �K�[go[�v�t�D=��#������_u� ;(7��>[�Lݕ4����v����!t�P��3_H3��S�²{���c-X��'"1h��!"&wE��)�5��D�L|��HnF#Pk�lĴ�J�"(/ZDo:�qa�I5� ���Ur������ch[K�^X�k�A�#*�)���	56�Y	���1�b�wl@*&�[��:�J�R�su��%P�tt��Z��Gmen�,"�4Յ�+*g����eӵ;�d�l������E-���1p�m�F�d��Ͷb�K�@����à�ZM��[��j�:��fV��EnɢU�Cm	Di��-ؓ#�+R�KL���[�tԚ<�p:�i����`�̠��±��L�8G:Ƞ���Gl�.�cE�J!E��fʦ�[���sp[B
����ʷ��[��/j�+ccM̳.��r�k�Q2�e$x���[FZ�e�f����سl�E�;L��l
��u1�t^Z)�����2�I�MZ&���� R:X�D�[ �#�6��۬an�4�cA��a6y�5��豭hU0��@�.)[mf���k�bBYF��-f��ф�g�֮�&`hmW3P�P9�P���`lk�W!r1�:H�&�b��^�X��q�͑uGeti	Z�m��M3%.��ִꌣ]l�X�4�"�К����aK�M���0���貔��t�6�)2����+�vi���\]3����d�h��y�Av�P�KYQÒ��fd��Rkb�j�G$ns���J�������l�7�wX,s�r��Y��MKn�8R�ؚ�&�@k]C�l��h<�9H64��昲��F���+���$.��Ƙ���Q�bg)���@��*�K���ev�SMXR�9�Ά��c�����&��U���kz�hj�rJ4ڸF�/:a7n��0���Xh0�1�Pkz�yMb\J=����U��.�eԀ҅���Gq�o3E�팺�M�fkh��ɞ���A+h���`9��<���㶆#5����Z&��6X]�H���q�$���?�ٷ,t��.���zX����uI�7��ʌaÚ����/WT��F�rZ� ]��7�*O<
�n,F�g)��%Ў��#7��֕È.Ϻf�7��g�.#a���><;k�b%��L*�T^z�\���pΨ�ɾ9�nꉤ�v��NON�lvG?M��(��z���l������1������Z�����Z:`�ۂw�.Ժ~s)�E(���f��,�ј�E��&or���%�Se�coμ��VwЦ�J؋�1�<�8���0*obK�&M�]����%��N�,�'����MR5S�@�m����e�+�3DY��T�L��9���1Mr4;$�28�/�χ��f|x�^���7>$u�W�;�uOHg�����).��:�>�z»x��l[Qyq-^�̧�X�u�v��_f<��j�3�)�����/�S��b�rp[�Nfe��d���I�a��رr���El���(�����rz!�Y��}�h�t�=�y)#2��=�dL;9'+\=B�iN(30e6#(n�>r���P"�;���r�u�X�=q3/�V'6����⃻�E��l�Fu�K�Ƭ�9���j�=�y��0;�w�C��!�.��5s�{<&��nǭ.��5�4�8Q��Bo�o���/LJU��[u!۟btPJ���?z"�G��P�Je~{��[[˥��7W>��3(��c�U�зPn[t��(]�kښ񨒝�&e�q����j�J�6V:��R�!c6r�YI[�b�q"A��Z�f�q6Պ�h�JЬl��u��Cv���W�E��E�,qL�+4i4���Ým�K��5&GF��-j^k5̮���le��h�	k�J٫����SV���i�v�\*��J�CA��)���6Gb=�^N�jj$*3�m�z{0�U��4(wՓ��%	�O'1Ph(�"�k����.�`��w|��9����a�E	B����,e����F���g1cN5Aݯﻥ����L���(Pp�ry��@�,&h�w]d�߼�I� r�=+�b��ʔt{�a5�.��Z�:�<|,�^M���K���G���mWK#�-�w�-)8Q��c��v8�>!@�ī�s���R�E
\�xQ�|:�i~��=�+�F�R�.��ں�2�d��ޫ�bTp��lJr�����;��5턚�_��f�K9��'/]���̺�VXu�ꄹIt�b��~�!g��T��K>)����&p6̣(������/V���-����2����&�Y�Ǻ��_�Ο[�%�Ϛ%�!0��jF;V��<ShM(��6u��ݯ)U�,`{�gpI*7�[/���l���%�ۈ�\�ª�ƑGo��q�Ds�*�)�bHx_(Os�$��̞$�IA��Q(S9p��3���H#:�ǖ�܍Ȉ��goj��8}�IY���Љ�#gp�#pǪ��YeT�K���S�അ�u�-����x$��ܾ�t,F�f�@&Jtč2od
����h������@�e�K;.��hV3����H ix��s@#�-�P� N�ZsڢT|(K�x���`M6T�:�5S�t��m��&�����s�C��l(R<=��K�U��(�¶�	�Qq���:�6�L��Wi5����H3��ۼv���)ݬw�K�_�g��fMw6!R��������,�^�
R��V殠֤�B���%�P�IH�7wz�
#3�͛JΊǞ�;(�d��o��Z�D� 67T�8�Q⒦�� ���"J��kw8��c,�b���p����Ќ�!Dȯ���Y����d
qE�v*����9i���-(��e��^�%ε�
�'aÕ-�f�#���+�����/�8l�5�Ҏy��9��'��~���~5$���I	/�>[��R�>�|�b��/�@���2t�&�h��]D���.���(S��̝�˹���,Sc�����n��滏�~��E�1��kf�}Ҷ10�Wvٺm桫�#ՙ	�ڣ�GC��G4f���Ӄ�����8ӏև�?ly�A�x1���Fz-�������LЛ2�j١N����ᛗ7w�xz��Q��j�����t݁�4�t/�H�a�$�3Sk>vO���Qȋ"���:����p�����"��/>��o�p隔5�B���O����ӝ�fh�n�V>�gz�&h�5� fH
�X�1%=��F�)���::.��G<����A�+L;+��X�[.�s��%��m�#�B�].�5�X��orw}��Y�Db����T����?u��A�����^fN�B���TA(��I�:-ݿ���_)0��c�M�N q�[R����6�5$�(�|2>99���`�w�ͫ�xg�o*�*�l(�J��ƢM�}MUK���:D��������߱�SK������^�I�%�mDa#�oKJ��Ϛ���|0���<s����Cd�R��:l(!%�%�Y��w��o)WA'Mmy�;q��vD�=�F����1������dZ3���K1��eק{gz� gzmKݵu�8�δ:!�RN�B���	�e	�99Z�mn�!�s{��<#�4�u`v�T�r��b�"�z�z���t�uK<��>��g��<��.��q�p{D�W��=o$�t��| ��t��]1G�ۓsޞF!�$&fR�(��}O���/b!�DP>�ٵ�	O�x��{���%�<Q�S�nJ�M-����i�I���h�ͭ�&˩�qg��0|�f8��ބ�4���,�R�j��)0��_�\`���^�ɵ����וg�CP�B�>B����4����ғ�[@�2�B�,�}]�9��z�� h�9]�&�%���9��O|py���FG���\�ϐM	�%2�9S5J���/����rjC6m�t�;��/D�|	�q��kJ��*}�^;M��zm�:tӨ!��߈^�P�P�)2�yE�Tx���\`����^U�$wTCP��.��f�f�o@"��
f@�B������̛Xp��0�q	H��Z�J9ф�ﾹ� q��qK`#���;>���/�Z��gw�v9MF���(��0��ę�I�}+�	����c��l��v	�j�fd�t�a�c�W�����9�#m�SZ��&�P؉hhGeD��ō-��c5ط��/{�Mf��aS�F�ٰ�]BSf�Y����1�A�k��`�Ud�G����4�vY�#���5Zu�#��l- t�Q�Ҫ�m��T5؛�f��E���d��%b�BٳP[,��+)r�LÌ#K`޸eãRMRF=��nX�n�۴l�2&�o�Ɖ��z>�MQ���;�˅�MV�������D�b���k �j��=��q�:jЋ������1�Ѷ���j��y[`fRͨ��[NYM�i5�B��I�X���t����{�7�C<��ͥ����w�e�ĸa�3�~(��W�c�?!H�bP�8a�no�ɵ��#�yK z���2ӧU*�I�Yܮe_�j�q	3�c��޻5�u��U��.3�"�V����xl$% ������3UT"h�9���Ã�{]�'K/��}<X��b��B�s����h�Yy���6|ʘ�ǆ2(10�P���E�I��æ�}Ii&*�o���s�/�jQKHHA
���iQ��<��P! fTPdId	�a2����	Z�d+fs�9Ήf�uy7�j�C�̵�a$���ϸڒiQH]a�u�h:P�@�Ή���u�W���@[���j���.����h�n[�щ<Owx�t�S���R.���v�RS
#N%��e�(�p�Ak]9D̦�IS>��4�v�P�1���v�&Yg��N<VF�Yf�a"hc��"�*;'��F�R�6&�3��q�p�����<�tK���2�MC?l�b��C���C�D�+��s����=ql�[{�u�x{jPx�I����
a�{O��X˪���,m� �8��<1YXo���>$ �H��{
:h���P� ����qπ�x{�G��W�YGa�L�������\�?C)���aF�"/M˾��,)��;�t���0r�*�rS�����&j�i,���7�{�vh��5U����r9�<�):s5(��W�~wY�LϿ�`��-[-3>�{��L�N���Jȅ�5V
L,6s��iD,M��D7������ Q�D��Z�!�pj#x!����ٮkdP��+Pdp��t��H$�O�&-�c��;߯��'�~���ϋ�'NN{)��O	OgʫR�B�C��"�k�kM�q����P����F�������\f�i$���y�ɽ(����ٮ�Qӈ���w�'"QD(�Ϗ{m�*�:4�S���$A�}���'H��|k\{<>���)���'	V5b��M��`*�h3��N�(K�Gj�*@�khk�U�	��R�FgW]/��f\��8A�m��JOui�De!�%�x�U7d�xƈ�$�緑�����t�!.�ѹ �!Y���v��ɾ����>�'�3:(I�/��K�2������8,ϟݟ�l̵�ٞ�g��[��2t	��=U���f�]ƀ���MtR,�e�(j�+؊�fy���Z%|P���N�%��u��/¿?=��q�E�������O5�ʼ,�p�s����I�a%9��Mj[�"������i�/f9 B�#F��4�P�s�M�42����p��f��`L)S@"��R�}qC�\7 u�Q�(�\+��/b�` �q�[��X*<Yο����)%�UR��YF�mwz�v�(��B@��[�״r'.�=*�w�t�F��$�F
Fi��#��7UCC
�*�*0\w]xK���;�5��DJ_
�S���4����=�k�B�=H��	��H��{b� �C9u��)0�Ǽ�X��gé��?xn}���&~Q�ٛ� A�̴��t���L�$��p`W>&�(KQ봗�:�ʱ<y�}~5�9\cX+Q�]f�ಏ�S�k\�bV/�L���G��Y�5�
sZ�s�G���$:�1�C�.���/sf�Bj�3D�Ob��%ģ��pn�mvY���Β� b�SuY��=��_V6�Hr�wD\���#"�!(wC���j�\5z@���3\l��9��w�h�n�x����T|$����l	�s.�M���3��y��_
K��вcJ�4T����@F�?,�=_8)R>RB���ӵ⏌"�u�E���*g��c_��O�� �6wσϯm-$�b�4<�L�R�i�&�hq���T�JY�{�"ӓ}�R}&��v����9��xl(�B��7Aj~�edMQUT_HX}����欓���Tٳ�����i�go���%Gۛ�8/}>�`)�����UQĨ�5%*!p��뵺��:{��V�I�u�*@f��>O|��8x��*��HӚN����aG�|��.��x/�,���tٌ}�@Ie������ |=��_h�YAۘ�~��^�)O��U�Yf���Z���g>j8Y����j�O��9u03O���|������L��&,G<�۳rs��Xq���k�+[�c��f�a
��E[aB͞L�f{]m[[��v
�������uu�f��K���
��5�kc`��m�*U�f�ꚤ��XXS�5���6���e�6�X7�ň��\f�RSM�G�ߺ�x�Pn
6�^mPT�ѷ4%e��X�%F�U�6K���k�)[�_ӧ�}���jѢ�bۜf�/v�����6sR��۾-Ђ��_b����N�s�cyNH����̶����]�D@��b��Ř��4�����Z@
�*[�g��3k*�j�����HH���F���(�@f�w\.���}�뒭�B��!Gm��>��rn�_K����i9u5D���ߊ�c���{aD�B�'�n��kNq�+y�/xg������ȹ��j]PܓEUS�}9��F�ŗ�ʼ��	"4�K�_�i�͵��=�;I�8n/Z	��5-�T杬,�� J��_,�qQ�\���5��]��{a$�B�5��n��}��a���TH�j��_K���2o	�z�%$��[��'�77y6�Q>iS��>rp\6"/�pm5$̘�:�@�a�H��v�-��:�����G.K#l-���F$�t��o�!�)��uJ�	#{6�7�p�c��\xg��r��ꄚ��Z\��߸.(�6{I
��2�Q
Q�C6`�O��xv��YR���lY�G�v�����h݈����9>x@�o��Z�&q}v��35#�����+U��ۣ1�B�j�;��}�T���F���
��9PC2�Z�,I�V�%��$F='�]�@��7�%$����G,���o6$��#Ԧmm����1�%YF��dY���L��Y�X-JbQG�/�d�^�4�n�s76�7�K�vC��W�ĸy{3�w�b�L����K7w9V���]U�1K-4L�%Ժ.���l(~!B���x%��;M�\�Ӄ�3.>?]Ԣ�p[�﫼���E|�dĕ�&W<X�pj��.>(��{�[<ͩ����8����|,�ɿaxB���;����}цe��Kruc��,b��fe��c\f��B$2��~���'�u1*�SS'4Re;6���ć΅_z����H��fvo9��Ti�:-<\�=V�^2%o�y%QRRi˚v���R��߼��Y��Wf��/�֫L�{����{RN+$�V�`=�k�$�P`�J���ϘZB#M���h-?n&��1�?B�F�*�^�#&��J,l�F�L�C��0{��	8��ʽ�e���]��RwjW���(���5׳�lH�b%�"71�4l-�B#j1��2My_g������������q�ˬV�q��w��s��m�;��{#7������f�,�K���6���e�X1-M
����^N�׎�,T
���T��s�=�rr�N�LL�!�:��Nm��
�iB�L���.E�ڎ������i�p�0�rه��[�g��uL�Hoy���5y�Q�{krgM�x<-
���B��[U�9�:��j�����c��#����*ꑴa{�2�D�n�8�i%�@�{.�<�&%��xo�?oz�ｋ�4�S�Ʋ
� ��𑲆uX���}ݽ�<��z��O,���<�N�`}/j�y>w<~�^��5�	/I7Mb�Yt�l��Z�S��|��E?[����E�=�j� 8u[T9��w^�ݾ�����W��ގ���A�kA��~��n�wW|4RtY�J�4g��EkuU�XQ��8[cq.b�1׹�C	�!B���}C�,5�|�ݯcv���g��u�zi`ѓNn�wk.b\s��w2��E��y��vu:YӅ��pLD'r:e���ޓIwt�Wz�}>�ǟw����2eF(F�'ҟX�=9���� ��K��Ob�lB��(��뻷�V�)�X��1Nb[�V�a�N�˜q3��z)^�zq}{;��L'�O���IG�k�Q���NI�eY:F�N�H^�}nu��>�ü�,L�.��T>��c�Ӄ&8�'LNme�(i��v\��T��1]�
�"')؇�$�aaٳ���Z�K��Pp�-��n����{��ݶ��sH� �;�`k7ߧ{m]���0�c{��5��ݗ�� �,E���
>|�����W��#��.T�eW�M�LV-*�b�h�t�#�Hl��B�,X~��!/��E/=�����ˎo S�ʒ���c��Ƽ�:W+�܀�T�W����vM9�m��nb�^Ѿ�6��q�*1Չs�ju���ܡV�b���+LZ;m��5v�o�:ֵU�ܓ�(OdgnE��.���{Q/oŹ�����N6��|h��ǽ���a�q�+�~Sw}eN�J�l���J���&�4F��j7�WsY��ٴ0N����������Ȏ<'�BFr������F6�^չD�@���13�7r��A��uż(�طtz����}q
PDԞ�3�(:�������p__#ڔ�ץ?�3���{�͝��;o/*�x��z��VH��Q]��0��{�I_v��$L�C��E&���*)bWo��r��T�7\��ؖ^ԉw���1�y}�t�a�P�t^oL�܇�"�%�Ϫ���]-�l��W�!��A�ؽd�����T��U^k3{{j�Cو!r
g���-�F0Χ�j�۪s�Gf�vs˱U�{��t��0�2�LɎ���ǗUj��[A�pF�����ݙ{���n�Qr��D�'������>M�t{���{U���N��/Ct%���U���c�-�dd��Y��n��6�����ޙr�}��0O~��I��ӌEl�*���STL��&�:.z��V�DW �K�r̺Zï������p���. ���*�����$��١� oWQ���t��|�r}��CrT��^�Ǳp�a�oh�]8l��҅���Ӎ�(�%"��7w����a�g>TU ��4�5V�,y��k	�MlDJ���ɧ����>/�|z�N��³������{��%XglG�Ú�k�Xۦ�ns�]�Q\�C[t�Rن���;ݝ/�׫�BM\�)LJ�q�������PùR�����[����;�Ԕ�J��p�y�3Y�k��K�x���2��È��ӎ�j�DB�6m�±��Ix������_��݅�J#� J̮/�D�3RI j�
[)��[V�-��M�����0�H3��	��p�m�H��Cܳ��� R�U9���+;=�QI%� ���q��xY�{ܬUW�	:��Zd�q�𙫋�V�ϯ]�l
�QQ	��=��)������I&�f��Y�Q�u���5wvUf�\�1�_ȴ�r�5fl2.t�pK�N�TqfK�;~~�������Y�����l����Ն�37-7�P+�Z�����gm��I'���Y���sjp[U[�`�<�)nEgˏK�e)m4�9�v���YY����\�5(�J9�n�薟��x�8��������~�2-t)M0ƨ�,u�8�Vٗj^KM���2�k��d�
��x�%�yL�R��i�s�$�ߟ�k���.��*:X�>�U�~DJP�0��+�N�Ϭ�f4�RS���/�^(��6����	��%�:(~���[�p�y���n�3��ޣ�8i�bsB���J\Ӵ��Ǿ��XQ�,��w��	
!x_��_/'�a��+'�dS]�3B�eB)@q��0������_EgC;���8z}�U�\w簑���j���<$zU��*���MK���D����~��͈T���#o�u���sn<*<X�o1^%f�?}�2dO>n�&��8�z�k$u@{�kB�,�T����P���M�;�#A󼒣p��FDb�]0!����E�ӳ�� �����߄����.�f���嵃.��g4Ύa)�ٗp:�[L���L [�	��چ1�t��k.Tob�X+�e�t�Ul�UhiT#Yj��K3 �ۄ���ʎ�bq�6ڈ���&�2�Z�f��5.��%��0��FP�It	t�B�HCS[��6��.mv�a�Z��%���:��9#nMpL�+�8+ġl��+L2Ƭ�,!���+�a1wMI��i	�佮�ZUJ��n?iy���rx!�l�ܳ���aS��r	�\��uۡ䞋��K�hF�J� �W�\�m�b7^py�G:���`Mձ?�I��t���=z��*݆k�͕��4�6c�tP�����l��#�@D��+3x�,>6��Z�-eAI̗�IӃ������Ip������//��.��K��b�m�����F�!(����s@��@�T�M:SC�>&ʖʣ'F�vi�I�,>�mo*�*<Y�߹q���S����X�I��߃�?��Hr���t���8�)�s@#��o��VY	+b%"Q�~�|8y
̼f�i��)��jji�	{I��/����D4�#��}>�%�0w���6@G݆��>x[��>}��꿀��ꔋ+.nu�ph�D"�-(A��v�jju�Y�a�ӠN��S�_#)��R�j wO}48��8|���G;�^Vq^jP�d-:f��G��.�.�	��'?xZtQ���d߀���'Dk��}:j6�9O��$j�0#�����MԘzayȥ�L<$h���X�	�oݫ�|8_-�>'�h\Ow[0�c(|�ϙ믹>.�Q��[''H�=$9��[����e���� Ƅ�0�T��4�D�Y�;c��zE���� ~a��z�����&�E���r���lBp��<0_�w*�өA.h�8�p��1^h�w�O��� g�؀�E�BŘ�Ő�v�ᩒME:t�!3J����6!JQ��%)��J|����ͬ(�*g�t���1!$u��g:_�Y���"�qMQN�r����\:X��̸�D��ת"aB��u^�%fW�k��
��㴨�Ø�R�,R@�4)�C�.Iu�mĤ��ݲ��
uk#��	�f&�
��$�zw���裠��[w(CFg������ᗍ���V�g]�Vg��� ��",���/����w��cH/LIqd
;������^=��g��a�<+/9~���0�J_�WOlD5�@p^�y��~sR�luTۚW�,>;�洋�f�v]יU{ތ=��/��E�wη#"^��\Y���>�'.$P>����
�K�b�=9A����w�y�U�U~\���'��������8rH4��vE�s'�츍C{E�{Tú�Ƚ|������p	���L:L���Jċ���ȋN�}�^�3�z(�Q���Lʁ��6X'a��I-MT�;�{��
N���qh��K�{e���p�r�_��jP$��n�^�����i�̅QUM��-,�b�V|_�ｱ
�\"#M�y��_���siQ�Ǟ�;XQ�.���e��Rԫ	w0�l#�mf�Qٔ���9�R�i�CX$��l��/!B�*��E@��P�$�*ݽV���W�Y��!�]������{��Y�\9�^�I�i˪�mL�s<�w3�����DY�|=�z�b$�4���_J>�^���jP�"'᳾τ-&I̲����)0��Ӣ^$�b��~W�ʪ؅P�>3ot�I�vN{�iQ���K=&�&�R��|�9n}�f�U��\���F������%	ï�ɭ>��zo��G}��>VT�S���ޕ�4��:���v�!.Ý��Le��Ea��o<ta����d���m��T%�	�dQ#у%}�3ң�/}s����ސf�oȋ���kg�<McDڱ�1�-f*s*#4��d���	ά��,��d�N@(�Fe	��F���-�L�4��'�BFg;V�+�+kK�����Vak	'�-I{�ĔP�!�&�����%)�eʹ�Ǯ�6RRB1�._ݞF�l�K����N����d�&ꛤ"huJ�_e�7���L�p�ɩg�⎔F4��_�zG��
_����ieOv'�DMA4�S���n�fe��V��!.�Iߵ�{���oXI�e��E���ȋI.�4����(R��
e:�Nf���f���`�4x��j(�  xi�0�j� �36�]$���$%�� �9�������߼= �����XG�r_M��J6h��� �5���x�?�a|H�Fl�e˖�D�ST�đӆz��$̏�������(qNt��e=wzX n�{�U>�eu�g�_k���2��g#+c�s~���,�#s�{b���~���>�ĕ��!}*�G��T	�ə�.:g�T=\C=<D�[�LԐ�)N�2E.ڄp� �m�ذԵ+s�-��Z��l��+�Cbl�Vԙ�L!1
�
f��V8kͺܝ��Kչ5[���.���s�.t՚kn�P�jd��)�S
��.t`m��V�Y��q�����R�6iB�Վ�h�m��<ê�2���P�5K�\\�Q��z��ԉa͕��b�Ne�͵QB�Y��{�}<uj��N��K�s�ّ4K�YM�. ��
�!��M��,��[�i�r�݃��O�]��]��v�/�,�2�R�Q�Ǡ`�"b�B��6�f��ΛY�f���Q	��L�cN��&�uU7�p���t4Dg>5[�<�W����#��Ox�3﫼���Exz¨��r�h��N�z�Y~�I�$��b�y���Bᾯ:�R|X�^�K"!�""���W�r_��2S&I�/�?�kq\��](�ײm)�	���fVlށH����6r���8�I	�fTJi��C!5�Q"��}[��|+3y�����؟s8���S��L$ģ�~���|�Y]r�朢����t�~[~�|>>��R�P�	6o�9<*2�x_�w+�\��$��b�X��9��*P�dKB�j
m7]6ͽe�1��4��-J��� ��*���j�ĉ�Y���z_��.��W��<p�s96saD�%�����q{σ!w'C�4�eEL�����(�>�Z_��lc��oN��R<<������=��&6�օvE�۩=�F�����"1�uk���T`6s:}��r):T<���
��q�����[�߲�[�{S$~!��>R��e�3�Q�diM7�tּ`Ё�rp<��F��þ�E
~�������p���}�J��Bw1��[
�B���Jf�6ɇ.���/�͛Q�a���kĕ��%$G���f���{�/�.�2i��$Ӣjds7�I�J%� �|ݔ�|��Y������s*���t�P�Q�D}���6n�ݶ�@���9�uSk
:C9Y~��vc�;�/'ú6�t���a�"�kﯗڞ��G��7�<�Ҫu"r���k�Q�,XAݭ���F��Fb-����z>oX%�(�B��m^��Z����%���˾�]��m�;����߬�mI)�QI���X�ΰ���g�O��&�Z��t��S�\-�}����[8:C�����&T�����U��,�R�������lߔ��l�� ��Ea+#���8�@��ĺ������D�#�S#	��#'U���;Ǉ#�o���F�&:ǽ�����w��V�.��%䗻f�-��)B��q��:q�� ���#r&��D;�Uw��}�>خ+8fI�酊_A� �2T()��ſ� �g�˧��գ�Yb�}K#��}�
ުGغ;upF#�DB�J �5�%������ /Q �ޣu�'��ׯ��J7�>ɪ���t�h
2hTPق�pʶ`vA�0	����쒖�8'㻣����e�DB^2���\�K�T�űП�
 ;[�=�O|,�(�2L$��j�u>��#�׽��/l�o�&2����p�q�f#1�-
]Q#T��V<���z.[]�>� ��d�:�gT,��TP�]9�0�)�����DCJ7�����N��oY��ӿxz��M�0g�9���b�8�jⷰ��������{��6fE'{z�3�3�&%Wjw$M%��q=��v:���2/���:̼��5"�´���^�o���˟���C��Ӝ�|���}���fsׂ��[=+�t�v{����Y�M�l.�v~����U8��f����2fP�ׇ��-˦>���xE�P.���{%�o�7�����Qx�V�.��6�,ғ���r�2cS�;B�������w`��a���v�Jk%���gvy���/+�\F������BZY��k~��>�SuM1:�*P�gl�s�[��Tz���~�Og}U2�%eVzs'.rg6B��� o4���'$B*"'��%��ggE���������\�M���g%������H���/j�}�
��}�8��_G�~幏��q��p�!.���}��qq���U"\�-����{�O�T[���k���t��mwsF9Qf��k,���w�	�3�_�h��J�[�2��Na�N��@
�;���C�廏��ͥ��:�=ہ�N���iR;�U{yTnKNZYxę���)ؘ;�J̲$ڷB��ПL�Ȝ��V��N�B��΍��ս�w���� 8��z�j��eŎ�B�|7Ӗq�wx�r�tc��lwOb�@��{��5�AI���ڟ���yR!���Nu���r.��ȍεb0nҙ���/0ܳ��UP��7l��[�J�9Qy2/��w{+@:�C�af�����(�s��տ>wI�E[��M�ޝ�%,�Q��Y���Y�̌�z�wU�'�_���&p��J�zx�� �A!�,p�>��}Vi�Oc���Ӕp�V�=��ORʎ�Tt";����EsLp�Zt9u�$DE#!�^v���/Y��&�R'�3:�SW˙�eF_h�aؽ\,B�B�t*3��E-��Y���E����t)�xT����t�+#_����˛�1������>g}�x�Q�)�I<V��-���$��2�'Fu���^u����,����Z���*�C������s;��ݠ�eϲ�q�	͙����U9k�4r)ӗ��Y'ֺ��H]���	3��e������;��숤g3k��Cmq��S��׏���{���,Y���u�����������<���\��{R��3��KT�W�/��k}􃲻y���B���ȯ)Fq�E�!����e���c,m1�E�t�ݢ
|�|q�U�qV!�{���O���zsR��6��eVO�ƿ���� ώ.MOb�zba���4�O��'V��z���Ok޻}U@%��nX�m��\�kVń����o�-��k.J�U��XD���^a*�Ka��;iQ�ʅ]]�&nuA�x�c�j�F,КfhA�Һd�bl�����&9ò��艬JAs�jZ�T�P��í���
�-�"p��e��U s��ٚZ`����3h���@�k(���-�6gMf�2��::[�2�.HT�&�Dĩy3��������v�hʬ�^�0�`�c�b�Q�Y�+���,y+H�Z��e�S�V6X-s��2�p�,�f�
��'T����mf�v��SFbБ�aZͨ�L֗�����!�!Lj�J-e�$�\$��鎕��ő���(�Ք�fp�Z�L�J1�x�a��g-4H��sŌ�;l�WG;]� Љm���m
�5h�)�J��U�s�čtn�M�-�C&F�21p�آ�����5�m�f������5���T�h��K�w���.�E���n�����xԶdvK�,A3i��ȱ�c��54�BlL $i��஻-��6M�̢*k�t��Ͻ}�2��4�l΁�/blJ�4f���S���l�+i
M��Q2�a��Z�e֘�0h���Y(�٠�])���4�U�e��2��3B�Z�{Cc�V�4�	��爓M�!p���1�K��ո��խ-���x�4��ð�5�5�YhZ8u�v-�P�,�[A���(:�hP����9�����fXA:�Q�%6����Ziq�u������fhҁ�Kbv�P�����`J�L�膩�Z�bdm�],6��Y���.�-�ޫlPi��)t9��^ٛC0c2���j�V��mK��g(d�N{`�(��]��sa�l��%�Z���n[M�X��3%N3����r�Q�!�N��it1(8p:�\���.4Z�K�B�͡2���Ŗ Z�<ڴ�H����TT�Ë+v�Aٖʻ�E!,r\*kf�mƔu������_�B��-�9iTm���{:��7^X���U�B[ݸn�����]��;�f�C��sN�K*��� �̒�%��dŃO�3�ދ��Ǻw�Md����@�%��'��0A�	(����)�6��W�����E����|ꐸ��������8�!,�v�-��:-�|��e���d��zƪ��nO`��{�쨃���Yc�{-����L]�:�1CD��Wj�u%	���[��lcU��=���?g�-��xt�M��4u	�>�z��t��|=�q�u�������B�����nz�xۓ���,�:�_�d}������iHPs��s�sq�bd��������-�y���v�}�;�o���\�p]�AK�{��w�^��d|�Gp�1�gʼJbV��Ƕ�����|��M���������u��z�87�ty��;�uZ{=�:���SBf���&�jW���x(K��ov��3=���Q��r�˵w���g+�U��^}�*C��Q�'k&4Ww=��QY��N�'c���m��*�����k�Lpu�r�W�rmlK���m��#���>у8��n��WF(!Nf޹����[K8L��ۙ�`�ai��TK��]j�6���;a��Vk旎�Okj.��)¥�Fg"�����Uu��u���^s�ʙ��6tٯ��h�K'i�>\�.>��R��yS�;�gb�x'z�`�c�%"Zj%k�u�l`��˥�a�zW[�1v��0��f ��Gu#�ї[��e%(�e�]�7mDۅ"�-۔KFFhɶa��̤�ă�.6B��]b�g�6��\��7�+f��j��n1cmBsJj�:�
+lf4����YR	
�.�2�����-Y�F��B�ev%LX�\ED��IGF�Xbgl�$�e�B<�FG��>��,�GE�����`d�܂�'�ˤo�{���|Nom�:����ws_�Y w�Q��8pj !�+p����f˫�nԠ�$h�,5归.i�ş��O�B�1i!2a�%=9������cO��x��	�iu}_UË��dD.�B�P&f%BGgDf� ,{·.G>�;�s��[;���鯽��Q�oD��BO�@�R$#	Oͦ��bvh��'�'�+�~s�i��Ͻ�o��%�1IMB()�K��������e��%��L���}����ϠU:Jp�'���A� �\���]����A>'��2SW�����w���{��
�6�Ӧ�R��[Q�,�X͌��Y�԰.��^�IP�)혺��,���-\��C�ST3[W�2w���MӍ�������{�]��r5سq
���MK)�n��߮{>�̈́�^>�y����a2�����-�{�	��^�?�ͳum�=�~z���?`utt�:/���u�}7������Ӝ4gﰹ�[r�k��ԑ�ղJb/'Q�1�ͥ�m[Dylǯ7�AɃ�gFuk�E���N�4$u5#ֺ$rc@���q�Q
�N��<����5�Ӻ�ֹ����n����G�@��!BIJ�!JP����qY��;G�<�$�}��};U���Nl���q�%�bL�����%��7~�����=]ϫ��x�؅� }�K�	t�2TLH��>�������n�<�����>�r�]D�q<���������w$aJK�[�s5��g��"!�e��q�C����0��w��k��=;00 �){˾7����d�l��]?{ޱ�gâ.�t��i��B�H��h��~}�YR�B򄰏���+w9��ܫ�������{ψ��F}}L��>^�3E:�~\����+���?b�2/�[��+H���G���#��ck}�s��w%�9��V3�q@�#��'C�=���3Asp���jf�'��W�&"�æG��>_SE��Po�������qmL�]�6C�d�?��FU߽�ڲ���#��p{�h��yߊ���Y���bW���˻mľ@���Q�& �3ѯ��}���񝡲����{��2<2}���=��}4�2hr�\��}��e}9���P�o35c������eq�us��
�Hz�@/����6����s7i�LcCm.�����e�b�
}\��r8)p"��sS��K��u�h�Ӻ������g�kT��Kn��50D$�H��<���շ��~ a��6�����]�u>���G��
~��I꩗2"�S4�_{=��]m�kv~� 3�q���y�'�=.��:�-L4T��}�!�RD}�O�};ȝ�#jܶ]ox��s�/=F��Q�4hu�D�+mW9�DU��i���E���=D2:�GG[����m+��꼜ܺM�Pә
	M#W�H��]�b�x2 ���2�J��N=�V�p�g�i���~g=���#��e��z����iX8���m&3����xc1q�<�"OE�ٙ���O�pDg�h,	%>�Ra%�{;�T������g��,[ܵOq���?�~9┄LH��$b�J�������+	�z����P�ڵ)�:O3��P30��2a%E���z�\����no����#��Ϲs����ܹ��:�hI��1)��&�~��x3�~��jT�h;S�&î��x���?	IL�"�Dʔ::�_.�n_K�{� ���|7'7��,����S)(�߼<ǽ잿��Z����1;�6w� �#�ߩ}�t�@���A���Hroa>�����x��G�f��������=M_�:���.D�E54����(l�Į��˽��ٶ� ^��G���C�~�%E�>�y �{�f��F�jÆhvGA�����ͩbn�6r�|�Y���)�n��ʕ2��D�K�&�r9q��^��U�RR+���Scm2Kx��%�-�ڐI�S�1���`�m���)4�)s��;E��J�ݚ[۬�Im
L���V6����0�1o1۴rS�3#��hS�5���Ps�����fX�m./P�G\�M�-F�KA0*幒�)	W�`��K,��e���(Ș�*U���Ɠ��Tq���
�)�����$���x������^�[�7��=콌�^Q�fj�\�rv� `#,ѻ��25�si#]�-��Id���Xl]�����*�����m!6�-DO $ #@ĐJ��/LJC���ka�t�.v�}#��h����'J�V�#��ADJF%;a��F�|<4z���'����{]}������ ||1�9�fD��䌣R���I���j�A�ݫP��x?{չ־���';�-C��T�D˨ngʻ�
R�}��Y?��m�R����������:oY��=PT�DJ�
J�:��pz;>��__��]�7���e������Ik�	��F)�)S`7j�$��2�n�´��E���M5���ϓ��*��B2���(0��6����^ַP�{�̽��Ȉ�>�ff��ݮ��^ԧS)0R��t���o�{y_��_Ey3_P����K�,w*zIHY��^���@#ԹV�6P�3'{0J�>��B ����OU��C�(�s�z��6���vu�O���"xw��]����e��ꆸ�dNށ���7����Y�c����}��	ѧ��֍��[WwY��R�!-�7*D����P��&�e�Bzrq7K�{�<<�������þ�x��+B$� ����b=�O�nc_C����Z���������ξ�C�EH�HT�L�?{)����^�K�!�W��B��F��}�|*6�O�Ǣ}�EL.�c�om����Ơ�(㍜��R�ղ�ˬ+��	MS���$�d�HuJ��;=5��/;LSv� g��Ξ�%М��4H��ʅJ�It���菽�޼��
�S��^����E� ��#�4�!�>q�(L�%c�%u}yܮs�n�VO��';Ә��B��B�c���!,5�1D�~q�B��țX�H�<l,��C9(�]0^�'����&r,���Q��<C3��N[�φL9�ߣ��`��u+��B��|��8V���}��`O*ҕ	aă�,���]�ک͛/��A������}g��ӎ�132�D�PTBCg~���z�.��T�O��t����w#��y�Ͻ��������BI�
J$�)(����u�5h��
��O�������N�)�C��� H�|"H�"(�P�Zء��t�X�'!ln���`�%�g��q6��$�hO��T��Rə�z���;[�;l9��X�\d�=����1J54:��1�3�P��1*
P�N>��a���r~�F����,遼�����nf�|LDr������%�N�F�/����G�x;2��wY2�.r���%�e#� DD�{O��^ L��!�#�T�����C߀��w�!-I���5�* ^ˈ���P�6GY�+�6+*j�_7a� �x���ۯ�Vi�����~�͂�*DI�5�O\	��ͦ<�}ƭ/&{:UsBB���晥ؒv�P�0H���]�_��9�R�2��A�
�����qv�"�E��y>θإV��$ͨ�L���roy�����L��ߏyӪ{�����X���RO��g��λp �1g3v&л�-�[�ݚ����(r�Nx֦]�wJ�|69���)��:}t����6v�[� ﯾ��nux�#U3N��g����[
�}��}U�nC�^���y��]�׬��M9�nZ��_׷��~����r!�	n�5z}R�qgy�y3Ɋ�"���][���n����r�w�^�~sհ�Г�n�[un��L�uJAQ	GV��F�ʙ�xo� �]1�5�����i�}ձ{��{���\wӲz����楬�O��%�����Aq��"�U��Gfw����"�,u5F2f��%����,�阞u)G����^|�e�}�Wd^4c\�9��!��B�b��j���$İ�i����y��,����K,�Z�BZ4Int�9Ҳ�M�:n�d���j�Գb9�0M�KB�[Mk5Y��)L��k��2b&��M���/^�BZ�	����R]��W#X0b�L�&P��V�X	h۫�%��
�,&�Z˱�l�L�srl<A �hC%:����W�>����<Ǔ���nd��5�9A7���P>!˗q	vv�����F�ٷ�4.��C��8vj�&�$�\�!��cF�bb�B �\,ҡw[��S+��I���&@%�y��۵o?��v�۸��V������ӧﾬCG��H�31!H1*R�|�\�w���x��~�I����}J�A�	�s�x���t��l�L�P�JV<��<��ѕ]� H�~��{�:�e��H������ĭ[����i�K��U���� �vC!���&T��Q2��H����r�6� Q���g��̞�;_{����{�t�=�nGI�@R%�9Q\�8F�;)t�]b�m��l��Y��1	�?���>��
@Ȅ�u���}u�]�s������P��?e�.~����;�̊S&�G�$�;��������}[\���5�0Lfsʬ9�Xm���\3�ziנ��u�˾Vս�	��q�w��q"�ԅ۲39>ܻ�{%���[b��sEp���@��~Ȼ����Prӈ/�Y��7qۯ�nl°��i�mZ��]��G��eH�P���1�0���G�=��S�|q�t�m�� �{�|.�/�A����$�j���V��vN�}�<Ű�j��_%�|�oT�Q���&$0��PS*&bR���=૯�蹝����bQ��d�bI1/V���^d��Q2���Pß����v>��xx.��p�}��۷���;E�(�C��ॱUQ̒�2Ѥ�$clCK+Ae�$��iJmD�k)j�wX�>*��HF�u�W�(��B�U��j��c؈�K�ݭ�w��W�ܲ�
a��a>�K+�x}�,����G��7��-���˯�B�'m�&Y�w~S5R�2JS2I�t~\v���UӖ��N+S'��J^WP�v�s1��fw�MVzA|���9�3�#�a�;4	�Zw�'��=��-�z�T39���A���g�Ӽw��g��w�%7)�@w(��{T��I���6w[��#m���o�-���ԋ��|z]"�5�uYƾ�b���I�LZ�ن��������2ȅ����O�hˁh�!w/o��,�,�w��\�Z�za����ۋ!�ʌ�5�sa�ff��p9m��*]�n�ˍx�n�ZBF����-�Wur˱�t'��MW�Zz������]�k����-��������Bh�����%:Mg�ܽV����^�Y�"�0�l����L�TȆ�.��tc���%����T�`�Q))�$�h*՛��l>o�-�Y�l+ʹ���ɆV��if�ّ1��>��t�2z�%��j�^{����w��U�3��I}S��������)q���{��wx�s@��̏�gkZd�^�:�P;y7�!���*���0Q�����}۔���u���6�fot�^/C�����e���	��ݣܨ���w��bgt��=5��.&���_���;[".{`��=,l�gf�P�G`�qW]�&:`�8:9
���r��k�6Y�u�r㘽O��y7w#��4{���L��<r�}�y��g��(q�;/�'XJ2��qD�"�lA���C�w\@�Եi\-[YƯ�ó.��ě�Lv��1^Ӝ�Df���ۋ���5tՃ:{[y�������c��u:l@�T�q27��G>@���w�-�$v��QG�����u*{�tnxb��}���xn�MՓN�>�'��ei�,l��,>)�B���Z�gڐq��j��
A{���7Xn{(��:�	q�Q+|F�e�R�VRb�z�9܇-��qB��T[&�B|�A[
 2�jV�+HV��������]E{A�VG�e=��o��<����Z�xwz�4n����3����tgAB��f�	�6���N��s���P/!ay��e�	M���ι^������ǳ���4��S������^�sH�/h�?Y�Ho�K{���;݆L�gX���Tfk꧛�����cc!m滓�ۖ��+��m�����f��ڝ�=0�X��9'��vݩ��9�sA%x� rٞ
�"�׬���1��9��
%5�ܱ�w��G%�y��0��/���=U��n`(�#���贎]I�$��[��{pn/V2�z���;Y�]꼔�9�G@l;Cpl��/2�e���dH"��Ǩ8����=.��S�5�V�I}��8XM����.���#M�ae�?V�u��,A�2���z}�O���`���{��f�����۶{�=_x�s���V	Y�~�����P�R8��f�˹=��U�]�2xP���^Z������hx/Fr�p��Pv��(�S�\5'�ف��Dm�B۾:���ԍ��Du�����Z��ܽ:r\�x�`5��N��d*��i<F.�/Ol��\��Uy������ ��3iW;�e��\�'�U}e�+ޏ�z��h���2ON^�w�	��%{l�
�AC�dMG�|ȝ*b#2�JW_����VVd�uBzch ��1SM����RX�|A���=9��]s����_M{T/(�}_f���ot��)u#��*z�n������ x�v'b��|v�h�{��O�=I-��r�t�3i��`�m��k���ZE����rЎ��,ͅ�����D� �X�M룗�{��w����6#�	^�)Nf�6��b�%N'4�EDDBQ��'��0{�l��~�tW:�nz�gk��Q�JD���R�z���XPeJ��ﻍ�.]Ժh?���G�xnu,��_|6��=
O��O$I(�\����������#'��EL=f����N�k�0�X��j�Ml`��в+](0C:E�����;�R�KR��\d�zT{$�2>��.x��>=2�ƝP�L�N곋qÛqG��!Q�iz�Y,�U�\:�89q�bã�1���-��4��V��ǡ��(P�lWӉ�BQ�L)q#`K��|?~�_}�5F�wZ���*��ml�>�}q�D|��bӅ����j�]���:>(����l�5�[Q˛s[�)��ǙbK2�lخ�c�w~Xye޺�OZ��;O��;�T��}���Un����z��@|��<��k�0�8�&QSQ"RGj3l�g_�x���._}i���NNԥۗ��6!�G�̇��
t��,u33O��u�^�nFV��z�~������+�f��]�|9S@�J�4�{���Bq�}�
��?��᷐��;q���J��M��N&-�wM7*l�������������#�I������w����w�Ue��{i�ϸ*?��>�6�+;Gޫ��=�&�Fw_��#b}�GCF��k[ ыI�3���/.
���{���3�C��F�ha�����ْ(��0�$��R8�u
�^a�Z�hQ�f����T��:�1�ԁ�� K��Kc6��\Fm�0k����F62nI�]�6��h\���]l�B4qR��R��Xhv#��d���
Z��j�%sJ<��RQ��!Mԛ�b�v�6R5�V
e����K�m���%���̐�c`�cb�1��gX�k��:��d�k���R�;�"��p~��%��}����W.��/x����\nnr�V��ر���7��,��N��Д��O~�x�~���1�I�v6�Yi��F"S3n[�Q�:�k.nk�R�����y|J��$̩����;;���V�ƾ���ވ��X����3�;E!���?P�Կ����� 
=�}��Q;��<6�;�j��4�gw�LD\()|�D��u.��gg1w/TFb�:^��G�{�fvή���C�*��d��ob;�{�[����ܨ�ݝk�m��h�&�W�v_Pc"eH���r����Kg�=`�׼�d����uMu�ٙߝ��Bյ�ۙs)�v�[���%�ڃ-EŁ��kM�`F�iV5�rt�ɯ��cG9>|�}�_�%���t�M�O���7��=�����Ą�����*%�;-�| p}��*����~��3�Sl|�:�Ni�ae�ǑƠ�e4���p[��W�PY�̭��y@]d�C�+��O��{5�&Z���^O�j,8$�z���Ŧe��}�)ݹݻ��E�V���"�����t@]�κ��(��0��b�üT���Ͻ=n�l�N�u-��:�������o_��3H�*&`�ICw[�9Q�]4٘?{�@�<����_쩣�dL�:%G�
���� �Ve��L�t�����<=� ˾�:n���d��JdL$�I*1����F>�� ��ح��������\�{}\��ogWj
�Х:k�XF�i��XmPms�LE�i�`5��R�s�9P��D(1"!%(I,=3��N��Ӂ���y֥p�{ve�ڵ��r����b�2�Nh��b�Wl"^)wkt:{�b��gi>\;��w�y���I��JJ$�a���կ�h��=��m.�@�;��_?��E����{#FG������������������\�<;�����/ǡ�����<3�ڳw6�'��b�	S0x
��\M�Aɿ}_�>;��6����{���KQ�a�����^��Z�p=Ep+�����H�nY��?^���ͯ�z���y��*����i���}�7�ڊi>��gm8ݕ�{�c�|��-h��$���1A���w�Ny��Nz���؅��g:Vf�Oo���>������yϫt��hM&+��hݚ�bX�Cb�a�`�J���J'g}�I������ͷsQ�ϗ}=�C���u�V��ʢ��o��!���8��<�A!iU
S�
�{x�������{�GGw�V�Ԯ����ˣ�����
~�y�ud�S��b;6̿�����|��r�����v����:+����?P`Zu3.f���}�
�J�/u{�<���GS�����c�g���o��«���ʲ����F��� �v�=AGv.�&�**<TD�j]%φ��>�Y��qj���ӑ�qۑo��Z/�Ւ�R�|�}s� P*��Ai݅D����͹�V<5~y���=�� ^
4����'ql�Փ���%*
�(�..�s��π����c�����uK�E��~����+��ʉ�n2�.&�tm�X��"b�.��5IV[����³<��̔L��4���'oXq��돇�~���ǝ��P�:Aw�A�D$�Uknf�n�������2��7}�ƍ��˼�	5
���n�k�蘚ALn��q�|�N\�u��@�_}S˛)����@ �pS�R��_��c������"�~�61ɟ����	�����]M}b�%A�FAI�_;����>�!�Su�l�k��ϗpu�����%d����y%���K�]~�@���0����a�M�nc�|UH�W76Q��Hw���B�QG�Q������ټ#���4�RQ�]�+0����m\v,9@��Pim�6!V�6�J�Z66f�+-56��Yl�4)�0�n�`�)LYm�qFX2�gh4�ԊH�au��F��X�K��u){k]�v����4WF#\�r1�1+��RW[���p�&K4�P҃i��v"L�h�$uؙD%�
,�p)5#L&5t:�jXF�$�M�R[�"�6��:�_gˏ��Ʋu�:Õ��>NږuÃ��D��wm��5W�+S��h�q��G�jgl���E~��^�t�12;k�¤!4�,k5�Յ�v��+���o9�~�sY$ǌ,e���D������}�*옭}����A}�r_C�;�2-|�IKi�����o�ﲹ^Ԓ؅"�׻Z�����xo���y}�Y�P�~(�HBT(�h��Y흇ܜvF� > o9��wv�]^S��UH���1�ֿ��=�ۖ)��5��ֈ�Q���I.�]�{<Y�;^�MKd�(���;;���n�Q��x���'j�+��������^b;���y<���H��)6��[2���%z��F(��@6�s+sle2�ܒxx#"%e$aJ�H?�;���փ��\;es]Ӵ>��>��s��9����$L�2�ѓ�up{އJ��22���:q�[�Fon���jy�'�uDK�P3v�ޯ+3y"1rQ.Ȃ<�����)ӊ<��Z�w]�:�����������϶N�Uk�6������{{Lv�&�qؔ䶯Q�m]�9k���9��4~�
��u2��G����;9��n�jzulQ��V�����m�r�;B�)$%J))�}�Q��'g�S\��{���;��ޭ�X՛�&fNB�"��n7� _/���#�"�m���z~�|6���Z�[U����iRh��ן=]w��������uj���]H�v��Zo�w�p>�e����fYi����kZT�cs���M�2�f�Qr"&ȴe&����9}~��m�w���������lDqB�=�ջ;�rs�{���PE��i��5�xz�>�ãGo��;^����-J��׵���YRPD̂�_ԇ�pɘ�7=�Lc�x1�7��ֳ���rv+)[P�_V9���K����英��Z�v�+�U�@�B���0J�[�*��X�:����#f��GSX���.�T��
�&�Vcg���bM��{.���o��H�6?K`�zQ�-�[���k	���ݬ���30mG,����5�C�|dJ�12�B��� ���c.��\��nf[����<�W�7f}�
W�RI.�������N-NT���D���ɺ�^w�o����oaG���g[!�b9N��,:�1,F��mu	j6'LF�nƺQ���g��w���^K���aJ�&bes/~��T��쭑��>µB]�/��j۝7�+�L���)�d�Ua���b�f����9�33-�bW��ɛ�T�nT����)ԥt��o}��_x�&����>�|:��|"R31�EL�������|=�w�bؓ�}���ӌＥu�]D}!C�e�D⪉��`n�ux#����1c*fo� �e��37b��Y&=l�eљG�?��ز�͐Ӌ�Z�F�� ��e�X���XU!�ޑ�E���r��R�j��wX�ew���&bDD�bTɄ�Ʈ�uѫ�x/{�}�asb�NT�u/�9	ߔ����H�Q�a`ًBlZ�.�P�M��u�m��:����-�L~;�`y��i�-�M*:{'��շ�����#'��g�:Q�j��'"
L(0����;��S����'�,}'��3�߾����K����Y{ÜT$�$&$�)�R��}��.55��LN| �x<���c:O8��Y�C3R���R*%K������a����m��r�?���]�pr���F"	�
N�]z�����}��q�nwU�ѽ�zw��ǯ]�z�ϟ�����?k�o�>�+���T���?9tʂ��?����g�3��˗���0Tt�UfHj�n:sW-��,I]�RW~��s�R�D�AI֔�튅�n`��s�H�II۷���.w����s�7��>�*H�!,hl�{��m�?�����;���ӟ�������߃�����5�f�>8}�?�y>~]��._o�~����|~/?�oʈ�����K\W������*��J��I���i�1�����nP�˴��}I��?�|���������U�����s�v~?�vr��r�/^'�y��/��n~��zW�y/���yxy^�S�}g��~~�>��u¹4�K51���a�1�MMhƌekSk&�����`̭h֦a���\Z֦�kU���Yki���2kV4kikSZ���Za��֍d�MikFj��YY�Z��3-h�-jcF�f,d�Y��kMd�Z�3Me��ՍZ�ֆ�֍b�[SZ��j֦4֍f�fMef�j�Vh֬��YkFjkV�i�Z��1cif����Z�X�ZƲc+XcSYmc�Yf���Yi����dƍe����,�2̳Me�f�YkV�k����e�L�Yc,�XkLэ�Yk&a�3Lj��fZ�5k&�c,ֱ�ce��3,jkX�X֖3��ƵcLj�1�h�Z�э3V3�Z�k2�kMk֬e�kƵ��ՍkZ�Z�ֵkLi�i�2���kV0֘�ֳY�k1��4ƚ�5i�li���5�3i�3����3Z�Zٍ6��c-l�̳Vi�f5��kcL�1�e��f��1���fi�i�k,kcY���Y�6��ֵ�����kX�cYk1���cY�c5�����kZcZ�4�1�i�Zֱ��Ƶ�k��f��i�ֱ�[3Zֵ��i�՚��f��33kfZ�1��f�ff�Z٘��5��k5�l�f����͚�Y�l�fk6�35��Y��c[[2�͛��31�X��Ʊ��l�Zͬi�l�Yf��֚�f�m5���j�l�̶��fͦ�Y�1�5�kM����j�5���1��lkVf�3k0�f�ͬմٵ��mml�l�٬l3Ki�f�,e�fL�͚�c3cL�m6fm[3-i��36�k[,�Y��i��ffl���ٙ�fkf֙���f3a��k[͙�e�l�f[6fmmffl٭m36�66m366�fll�Y����ٙ��5�fͬ͌ͭ���i�3fdڶ�m�Z�͖�kf�i��lڶ6#a�l���6l�����f��k3ffմml��6lƆѳem666��f͛[[5�i�ٳcb�m-�M���dmM���jflٱm6�ɳ5[V�lmlm-�cjڛ3-���V�ڶ\-���&͔�ڍ�f��m[Sbm[�fͫf�e�l6��Q����16���6�6��lFձ�6+bfm��Fձ�l�-��jlmV��6+j��a�lM�ca�[Vi33U�ڛL�ڭ��6�������[[@̳-�ٳ5mf��Ѵ���M�T�L�`ƫj̛-�ڶ6�YY�6mM�-��ѱ��ڍ�kb̦blڛS�Ve4�l[6L`�fj�l�4�`�ll[3�ɚ��e3)����ٱl�+��&�2��1�٦�-�%�̦���SMe6k-�Ս��M�ڲ�mk)�6�L-kj4acV�j�j�a��L-�&1�6�4����5M2�j�صe0��e���1�ͭ�F�����MYL5Lj6j�2e2ac)�)��ڴ�mZce�lei2�bɚ�blѪdŲ�j�d�hb�2�Ƀi�T�յX�������Z�SC+jєє�)�&Z�M&S&�+)����1��b�щ�&�M&Z�&�f��-SK)��he4j�2�5MZ�ZL�M&�SF�+)�I�)���)��dj��d���b���2�d�5i52��&�S&���`�ij��MMSK)����22�2�����-&VSS)�T��ur��a�ժd�5Z�&F���iahj�2�ML,�S)�����j�MSTɪjabaje4�ML�&S���Ŕ�e0�5M�&-SI��e54��S#E�I���i4�YYMFSC)�)��ɪd�j2�LLL,,�F���a�i2�L�MV�)�T�i5LL��)���,YM&�)����0e2�Y-&�T��i0��M���d��YMKI��4�M&F�)������42��ST���j�����i4��-VSCT�dah5MSI��e5L���j��L����jXZ�����j�Y�&&ST�YLMST��e1ZLMSCT��15L�S#)�e1Z�U������j�L�VU�d�M���eYL,��)�T�12�����j���)��i4�XZL����2ZL-S%���2Z��E��aj�4XZ��I���aj��,�ST��iZ�SKE����2�XZM#T�e22��&�T��aah��XZ����b��YM+T�e2�MKTҵLSI��MF�E��i4YM�&S#T�e0e4����j�Z�SJ��i2�YVSI�d��,��)���M&�����i5L����22�����5M&�R�he5X�LV���aj����T���j�VST�2��SE���0�LVST��b�L�ST��jZ�SI�ij��SE��e5L������h����Z-&��bi4��&���dj���T��5MSI�hai4��-�����aab�L������j�5MF�U��j�4����԰����T�i40�XZ�L���)�h�YL��,�kCMKX�b5�֣��5�Ʃ�,bl�i5��V0��Ɔ1c+YMb�2��֣Z��̌�cT���ikC��cU�&�Z��Fj3+Z�����S0f��f�dk5Li5�YV5Y�Ɔ�Z�kT֫X������V�5��,��Z�֣Z�ef��5����f��cSY���c+YL��L�cK4f�j���c��hfV�3�5��SZMi5���h�V�kU��bc+Z�ecK5kU����&�XɍL��Li3U�a��ef��5��-a��`֦0i�1cK��Z�Z��ƭj��X�h�dkei�̦2cicC6�Z3�5��,d֓L��Mb֫kKZ3U�5���j�3hc+ZY��1kU�Y�֫55�4kS1kK�w���,ֳ���`�_G��DUW�⾯���ݯϟ��Z������o'N3��m���w{<.�g�?��s��G��>3���;QU��?Aˇ���~-�6{��7�;���O)�Mv�'��K��������E�g��~c���]U_D�M1�}_��~gǿs�Cۃ�/��f���UW�DUW��m�h�xn���ҡJ�=?����~�-�fq��w������C�D��y�Q�]���e��_���>/n��n�N3'�qw&�?�pk����y>�K��:N�EUj���s�������o�}4EUg�����n�p~��?#�c�p��{���|i�C�U����ne��?^����O�Ʈo�~���h����:}?Q��8��ƿ�z�_:"������v}_���|����A���O�|O6���t�Wa�7?-u�۷�u��[��k�~��|Y�ߩ�����=;�?/������W9���x��m����|^>4EUf����l���}?t���G��x���w�f��>����]�'�?�~י�|���_d�R��G�����?C�]<S��T)_Y�w7��=��g��ӱ��.\3���������?S���ػ���PVI��Zh�����` ������Ͼ8                                      H"��UR$�!U ���EE)"E	UR��T��R�J�B*A �%$��Q*��I%)H���*(
Q$�P
"�)
R�%T@(*�@�$$R� *� P
 �
 E���J�yR	R(�� )��R� �:*���C:�;N���z�纽�Xu�{��jV7H�7��Zn��%����n�ǖS�whY�&y��Zk�w�UW��i�����V�9��UBT�()TH���(@ =�]�D�A�8��x: (�^}���PPO�()�A�ϻ���ރ��A���ޝ�s�w>�*��޻�k骯����G�j��t��#��]eIG��TR�=�$�	*�*�H�+� R��Ů�U*���yn�m3���Ö+��管����+O]^��\y֞��8�t/3G.�gWh˺6�ғyB�=��CT��9c�y���%D���T$�J���{:�X�2�N�����ny���������ʮ�t�jP������q$�sʥX��Cٔp+cR�n��j���J��(��*�J���TJ�����AwN<(�^<��V��LC׮��T�W �{ӭ5���n��5.�ͧK������kݷ�US�g�ּx�үL/yQT	QUB()U@ Tps���ǅJ�w�A�
Z�����^���K�����r%
�Q#�����'*�ʮ<���8*�yk�gkZޔ��� ��%%UJQI��L� 
.t���u�����u�;j�˝^�u��j��x��������՝��Xw����W����@w��*�go q<��uk��H@�� �PÍ�Rj�z�PFu�:���0w�s����v�n������"�����V���e+�N�os�8��Ū�PǐUR��/z�*D�� J�
 L@
�
㨣�n�4��� w��y3����<ͧ�v��I���v�93�7��Ǔ:DֻWr��4��T��i�=\X����{�D�J�AR�(+�R��+��g=�t5�%I�w;�:�^��K�ӳx�u�J�rgy�9s�z��+�[����绣+�Љ@s��B���                  ����Pd21����IJ�� 4ha��5QM��Pd21i�R�bJ� ��$�J� 
Q�m*�P 1&BM��!��)����z�Xf:���L�o�ߌ�� �
�����@v"�� �
�ނ�*�DVQS���g���˭�}=םu����?4۞m-ѣ;su�mV�����佤h#�Y{{e���@��R�y�����&��ܒy�9��v�1�8$
���%WVr3�*ܫ��Z��܎_ȩ.oK������z�O���q�7�%�^�q�z`��W[��7hɌsw�i���قQ =�G������K��}���<Z�q���*ʵ<��:��f�b�{��#{IV\�a ]Ý��맹#��P>�G\D8y>�i=_ds{�.k巎�~7q�FM|�DO8��{WEh�Ϧ������pW��&���y�L���������SXK�{s��l\Bt�ڢF	��e�u3�����ٯA|�޺zh����b�λ56�L>�݁ɩs�LɧmԒ}w��ti�xhR��K�o�5Z^k�`犙��N8�k�E��fh�U�"cp�D�M�4�Ѳ�Ȏ�F���.��_p�w#���GV�":n��T�Dw>��E�#U�np;n�8���G���b�΀��=0��=���f��څ����U�;sF*�1WgA��==T%�r�:�m翌�^t�7^l;o�d	�e�I�b�Osm�w���s��7�5v��h�MFѸ�����ϖp�<��K(a@f�� C����<Ry1gu-�y�v��נ����:8 �\}��'�3
�n�忻ՆM4���z; �k\!;�%e&���GI�̩��7e�ށ��}�nl�S�nL��E�Gw~�����$�@Y�-�)��g5�,!������8�W��_(tX����l�8�o��?YN�`��%���7�C2��W�os�����سP(�g��o�`h���G\"�L$���3����A_r������a��[ݜ�ر�x�[���9tf�;{77nꢝ�����[��xӢ�3��9'�&U -�X�K��ٺ܉��4Dvީ�5�2
֩�6�1�t?��.�x�in�GF�N���Nl���I�.P� pn`�A���k]�c(�x��Jf�.W����;G��Y5����Wu�e�o��	�w��F�;�8Uy��s9��>1T�ڹ;��a�ŝlC[Α�����omHg`!�3�:�9�������3q5敶n��F��/m�0����������X�k�����F�C���;�"���&��}��\���7���6����0��7zN�&�,˨\PS�{�~ݡ-�A��\�tL�H�7�J�ئ5�U��/3�gM����9�J�q�0�`?�b���(Y�d�q\���9��]{�Hאs� ����4>�	B��[N^-�v�Z�;%U�E�	��^7�/;D�*3MO7�Yjk=î�d�ڑ0��N�po��Dm}=��2YFhVZ�z����ì�U����4�F\V��ްCVu�� ��~y�	�����$\�:^q�"a]}ݡ%vvKw;'1r[��:�Tl\ԉ��W<��&v��[V�ίZ�x� ��E�'>v	T�X���Ð��reS��"3V�=S����6�Mn҃N�Hk�ݻ:]]RR�^�+�9���.�I��R@��&�a��Oz�4�R�X��4���i���zwwqy�Ԏ�V�A[���s�$s��@3^��r���>���f��^� �Nqe=��2�l�,�Q��ѯ��8qmBضlɇz����v�� ƀ�zB��9�z�"Y�����q�x�9/�������ӷ!k;wk���!(HN%�Qt�,�e�O\�*;��Z^>�����,��gs V����$�]Z�E�����1s u�3B�(�;��_��9�[�� �J�%'�taʥa��\�V]Rtt5�j�&�:r-5w~Zѹé�!3��x��W�3�f�o":�Inܙ����mP�tv�Ferou��e�:��Ξ����ۣ��bԺ�n���r�����wv�
�xE�x�=��$�+pG�Sݪ7M�3�ۃj+(yqbjʑX{\�{};�z�l�sM�%�Bbc=u��s�R!vb*�/ [��od^��Qg7;p���bͦN��t�J�;��/�ӰNf�g����/&�ĤJ��;�Λ��c���*��@Z\�jP�=nwA����؄�	��:
�S���Ś�&mǺ�5�8�<$��Ó\������w�k͒��%b�ٌ� ��[Ma�ZU-��|F�Ϸ�z�G.	5����s������k��z�f���Wa�Uk;��u�L�n�r��2��iU� ��n�Z�=M��d����{����;@���f�e×)��%ӎT���^��a[�0������Il�? N]�4�WC���7r��'��6����Z�=ǆ=Dq�~h
�A�,�n�ܯ翁1)�������L>n�fqD�lgz�c ���p��n�允���Hw$�� �\ќ�ڭZZo��gq㽓6C�2��I��U�\���A�1%2.�Ӝ�6M��~���sB�{�WZ����=�����ɔ.����]j��5��N[��r�<��ac�{;
��sui�8:��r~ݗE��w)���i�C����W����k�4^f���4����m}M��[�-�͛�=N�m޵�ge���l'm�N[@�u�$.�m�o�u0�|c��و�ۻ5�^��)W�/5e�p�r�Qf�Ӊ��;���Y������Z�=��j�7�`�C|T�t��K��T��k]i:Vvh�޸�s����P������p�Y�ѦC�8i�Ϙ�����{V>�h������8D�<#J�x�����^K�&nCH����bDDg^���h�i��yQbǡ�'I���ȫ��aW*}Y��ڦ���Nwq�������x�(�x�m]�I�r�;��:�tn��~Jm���^��@qS��*������4�bHvP�4���k9j�%�8���9�N6{F�;w�isyvL\��M;���˿��)�]�qD��{���%Pޣ��&�F��mx�w
p�ꙩ���},��F���8��3Nw<P�O-i׫��6�fvl��u]��Ю�l,���ږ��=�j-�˿����CVr�k���0,6v����3���&]�&�0>�cyc`͋!zɼ�'u7��6U9�9�>�"z惛��;�X����@L�\-@騺]/5gg%���c�'�T�cc��\�{D��S�fn�7X�:�+\rԉι���m�I���Z�ő�ẓg�0:��f��ݸG�w��iK�:cJot�0��P�<�t2j�3�K�v��Q�p�y���^w�[8�rJ1~c�<h� �vk����~Z;&i�}|�k�&���E�"z�E�+8�ۚ�y���b�ø�RM�XǱ�8�R�{Nu�)C�n��mGR���I��ܛ3s��
����p-t݅u	q�JB�����M|�4�FwH�ͷ�aT��e��.� ؜3e�Y�� :2���A&��jR�C��������0�qlf��NCY���	�{G]���c��9�kn#H�0t��p�L�j[2f��j��$�X�ٮ�uWp�����;�͜�=V�����m�|
�w4�4G��1�NR^᣿�ܝ��br;��W�iӤ���Ӌ�2흄�z �n.��l޶Y�fB[�9s�r�ْw;KΤJ��}(�۷��iE �g3pR�	iL�'iNg'Y��=-�p4{oQ���(&�Q��L;��C��A�u=�"��'6�>|3p~W�=E� �g.�]<)� z��i[چ�ӓ7V��t䙹mO=��9
�?t��%|�R��Zw������k�8���Ghʒ�Ե0^R�tYuK�S���La`{�P�.�=�:���]ق �&ہ=7�ƛw��h�w�#���n\��{D6�5˜��ui��5-�I�v<��on�IYڰ~{�K�LAW�S�i�r�2�v9�͞#�(h[���V�n ��t�ԁ���t3��pt���ՇLɲMT�5r��RGaO1���Fo����5���d+C���җ���]#IΎe�Iu �����gI��uAWsJ�Af�2��Z5�.m���6e�h��B��M꜇��ܓF�1T�_���t��[��DG�����Ū!;1��x�Os��b�t��ܔ�ˌ��owwIѫ�n���Gc׃�u���.�p�J��e��+;hש���ê����k%~��{�X�z�<�͘�_�{�[{���o�r�ɂ�.	N��ػ췯#�h����yќn�ǀ���ӻi���n��돂�ь����ĮmbwD��?��;dӋ�[8��L����*�1|���{_,�����i����� ��?^ţ	�yέ���D�յ�G9���+N��{Aɺ7��\�8�q�f�u����I�5B��'r�M��ڠ@Nչb��a���pOj�����XP�W~����{��R"���n�M�e���]{7'���o���Y҆y\;{t}.�Mu��P�����y���
]p�nG���cE�b�|ι��qMZQ=��D�J��ٝ�ǅ�Ҷ�d��h��|v��"�^;�pOf��m�.wN�7_��ئ��5EMT�k��/=�X�oe�N�v�ы9�m���p<�`��(�h��ꙋ�7�S1��"�7�F���E���wR�
Տ$�K�^�\�x��9��5g$�����S��y�o���˜��^tΛ��ʮ�h]+�x�׮6�t�^޺{�eh�ĵ�`�'�`�zGd�N�u�>�*ٳ&�z��p$� �+���������AEhVݚ���I�Z�͎�w]�����!��]=�M�J��	t8�@�O��P�<��R��?��,��t�	�F���V�ѽZ�/��u��]���7��	+o�{r����	3O-�����Zz������u/7� h?m3[Uou��q�ޓr�r,VSSlw@un��;Z�%�y�"�jZ�[]Д�͉�TL�	BMO67ƴz��jL�_�%On����4GDvW�.�4��f�ڨN��u���ww�N���S]�"{���l�l�ue�L�	��B�ʦ��<����}�ou��H;�C��-���]k��o.@�;5���î����/\�����-KQ�8��4���_����ۘ.�������sN@\����M�JR�fZ������l#8�@bS�r(��Ǐ��2vn�@gZi�g`��=3U�Q�͍n���{R����"�����
'Y����WWj��
+�V�G;�6�u��,K��^?�.4U.��ʙ7t�Np�&1Ormf��N�5,�%�,��9Ցy�5��ʐ����͇�,���J����c�;�r��e�usݩ�1۱dsxF7P�܆0���?<&�WoI�N���+^��&]9ظ<;�~X�Aۂ��gn ޜk��P�d]�s�U1��ٗ��[�~�ѝw���-&�p��k��qZ�Ά�G��wk2*&9�BM�!�@��t��
�S�����R@JyT3��0@�`%�t�M�6���p��3��z7���h���wo�J�=�K����*�܆��V+�������HŴ0��W�&*��~]��E�)K2;WE�Y��{m^k9�e��Hp?�ࠚ�
4�p�w7�N[�4���is��ݨ!�J��t���v8�W"T��e��s�G�w!�M�V���hv���ً�9�YR�ܠ�#�腷�Z��܏fmݓ+Ԟy���(�B���k[��~�z#�L<w.[�ܜgW�[2SZ���;d�a'#�H����0ܙ�{�L�;��͏��n��9~�3V�7��{�3�If���Y��wx��]\u� ���Wo�:��Y���j~\\��S�Ba�.���,c.B�*���pВ��X�@kS��e�b��Q&�r�6p�{2�r�m����h�hs�v��f�+ݲm�ו�'>��.�H��[�Ӕ]���Q/�	#ͩc���5Hf���V8�8���Yy��Q띀C��rݼ�ggc�� ��a���h�q��(=w���U-�4�*�C�����P��n��zt�q�Fߍ�k�� �p.�9����1@"Y0�;qu���y��:;sc\��z�N���q��O�\Ѷd8��h�z�x.kú�gAp�쁬?��ԛL��� O��m]��qq��p]��S�1<�:k:C����JWxLٶ�a��[!G����w&�gZ��!Nي/�LƝ��"6�,p���'X�g> a�H���˶���j���sC�zk=��qe��r��`b��/&;A� ���ݯ�=�s���;1�e�u��HgD�7v�SR��˂e� X�ņ�Q���)���`����V�&��9��rw�Q#i���f�clbmw��Q�M30ڞЅ:i`G^���Y��	d���;;y��ܚc����ox�`�٣
ȴu���SB�vs�B+F�wc*��\��3�����׵�:���2�vK�ק�Yݐ��9l���z?��8ӛr��w	��z��#^�l�x0+ �zq/��0�ڹ3�c]F�E9Ű�c�M����K��A�Q+�($.m��h�P��4�6<x��Zט75ª�zp�on�#4IWmj�F��,��t;�i��a�g�.����1����ݱs8���MK5� �Z8��n^)e�s�]WL0�����DH�΋A��.�]1v�kDfd��a��Qx��<a�-��'1��A4��y��C���[��HR9M���]R�*�c�0@���%�a�[���iq8C@�P��?��:o9����Wn���&[kk���;j�t�M�U�gmP�\[��
Mu��VZ�cy��aE1a&��0���k�He�T��c��f%Y�8�	��]�%h�k�5��X�m�q���&�Q�ݖ�gm,��$f��,��	���8�����X��ʭ�Rd�RML�B�&�f�:��:���GL���U4!i	s��PH�Q&ˡ\��lD�J�����ɚ��q\k�6-`,�%���¹�����U��˕fՑ�L;Q�EM@���n2�:�Q�4ūb��,���h���j��:լՄ����Rk�!Ė����6��K�l�-i�d�gMcs�4��Gr�05q�����@hZ=�(܆���x��&λ5�b[L0+05!�Vl�SW8��찍�]h$�h`��[fm�K�[I�ۊ��c!V$^IJY��M�D#Y�%�	Y�ERԥ44�	�p��.���6t���Ziwf1CK(���V�	�Z,ɵ
,�H6/k�Vd��Z�t��0�v�e�D���+��$mX��Ӽ�ǆz�t�+H�f�f4KS�+-� ���	5�#7$���`�2%ֺ�Y�Yv(
�o���mW���m*

in.�6��ׯl��YY)]W��@��Es�F�I������mp���:){p,�Dk��n :]�˥tIuv�.���+�T�����.�a�i,��l

�ݥ��1@�lЕ�m�����L�en`sY��":K���[�ʖ�PZl��Q3�Ch#�e\�eͧ9�\�xˀ&)�Y�t�$20�T�l�.FԼ(��ڙ��*�
��ݜ%��e�)�m���]��R#2nL7VRbͮu�]M��eF�a.)r��(���(Cn9�̙�ehS���f�劄��ێ��T���
�:�	gT�f\�����(�ˎSP�M/f;3f8���m2G���-��mlۦ��F�L�"�&֊�+��S'�(���4m׆�%1b1�ce�ƻK2P�q17
T�R�n�6�	T�-�aũ5rZĐ�;�ּ(Af@��l&Hf盙��JK8�b8�-����]��k1"��m\M1c����ڑ��J�t��@�cQ0�Z�ad��Ӆ��J2�J�ܤ�.�	I��u��U3. :��2� lk����g�T�j�Rі����H�_cOhT�Mi4Ғ�e`	�H:�����o�%ҙ�1n.,���b	����j�a�l3mE����ХU-���ҹ�У���k�e�S��ƋY�5��k�Q�(MH���l�C[�R�R
;C5�&ʚkJ,��>�ɡ})���9�d1VXv�[��{:i�q�l%��g�i��o,5!�Ў�U63k�lF������iH�h�תM2c��G�b����6n��L �-�l�l��M�-���1�f-v�6Qc�]
��cf���-��y�s�� �u�X�Yp4�+9s���غL�co�oM�\��a�Q���d!�B�+1�[��Y,��s
�.Ѵ9
+���k��2&fmph �6;�H-����b���J��ӎ1�PM,��5�kod�j��э(�̚�����b�s�U��EX^	M�Mv��Є!��6��
Rf�`Y����j��Ƭ���mF�ˡ.��Df�[4mJƀ�`9eRY,&�!k�J��r꺐�p���m75�aM�Q��c2���=e��X�Yx�ڣ�e���A������s-�F�[)af-�Tai[��Y�2U\^3�贂!k[-_Ys�0Gf���p�[�ĕ�wZL����������3Z��.k�Z�-���jR�ֳF�ehm`��Ĕ���`�W%�����v1�Z�ԸX�K�s�/!������	�fX��:�KfNٖ3\�p͙l	B�pfƜ.ڰ�k˨[��R�u�� QG\�U���ބm-� ���m��4Ҏ�kM��r�(�bWd���͜�J@sYn�@�$�S\��DV3+�w-�@`����X��XX�f�2M�r]���a����l�	.��mub[]��J���B�L�i\ö��]�A	t��х3���Fa.��,�x]�����T�t��)I�G]&���dY�*;H+��
���ŘL���tc�MD+4.H6Ȕt�˫�j$Iuʨ6V��
� ���n���\�+�l��M(��ݭ)m�.u"��XYV��n̛1/0H6��7h��u55���bm�e��8\ˡ.-)�1i�J�#�.��ɐ����<�"V��Mp\:�)v�5*\^�M�.#D�]a��v/	��j�.XZ�&	�:�+��/l;�����M)B��22�;r�i�bd�l���]��M*%����1ĖV����P�\٪�&ű#��uʓk��4�P9�`��!4�<�"3Kq�jt6��*��<�Z����[n ���A��k{Wq&c��6� bdt��il-�Y�n��Y�ݒ��5Lr�A�Y��Ů�Q�ک3nx[x�.jی`j�M�ń/]r�i��;[�#h��׮,�s`F͛�īLP��Y:k� �0Q��6�&f�v�6jm	�n#+6Pb=kk,�X/8c��Ҷ<�GX[��B���J	��.�׆C��ز��F�f����=.�ae�nj�"9ݦ�c[��v[���n�6ƙ!K�^6���H�Fd5%m&�`��:�kMn��]\�`M�^ц��6���`W��[�L���n��ll�	��m�bf� t��#�e�֝P	�G5;p5���H�V;f(�l��h�d-v�\b⭢%�]��n���.(��E��2[-11Вڮ3 �4�K������*c$��rhҷ{h�c��!P6(���f��W��	h�`]���pm����K��&i07h�R�/	���k+a6� �H�1��[���[4�͡���"�f=M6Ҷ�e�&�W\�9�5�1٣�9�`�7##m�4-�.�����k��6�6ڻR���30���j�u�f(b�.f��]jWYIf@���-��#�\Cik��S�XA��P�̈́q�ar�J2����,n�XD�
J�[m!`0WPm�+*jVGVWJY����9Ġ�밌�#6�i���q��5�Llݝ��4KFf��MK� �P�ڄ����R&�!4�WFnWhՖ��&c�[�0���0�#6G0�nP�!Y-flR;jj3d\b��թ��Lf����[�t3K��Lmx���冲���ʰ����h��Dt)�"k�
]x.3��f�,+���,�GGR�R��)I��f����hSc	,��6W<X�����0����е��Ќ����6�Zq�Cs�[���4�7b�!˙{B��6��"�4�K�Y��Rע�^�D�[&nɥw$�م����\d83Gk��2�49q㵘,��c��W8捩�A�hg;v),q�[�,&��COx����u��� 3.+uXb��K[+��)	�6�	*l�Ƶ��m�ęl�%F+��h)�8ۛ�ڹSb�KT�L��Ym�N�2���E#S�B�c���WT���K�rBg-/ide��bgi��kM��m�V��8�M��J�-w�K��S2�\�Kp!5e��sb��A�0�m�Ε�j2���.��hŻ��XQ�J`V��iZbhi����Έf6�^��q��a��ΊGc���1��X�]5�b	K ����a����y�ʸ�#6�P8�pkb�F�+�4���u�Lւ6��ǖ����IlGj;�r�����X��c����kP@�"�]5����J�*��t��b(�[Y�!:�J��&�i���6�%I��6��V]Bb��ܼ`�-�­-&Y�Չ�G���N2%���6����/js�ېm�%�ؖ��]x��"P�@�5��u���2� M-p�@�f�؄K2�X�R���U�d3t���4n^Ժd����h�FfXj/4Eƣ��� Ħ)j@�C����:*D����Ia�o�A���3�@)c�&�es�dH̗P��I���������sc�,t�v��Dq����[4c��k���^9��u�+��8amJKδ�M,��5�d\r��m�&�f4%��A\v36��h�VU�t�MB�CX�k�����bf�+e��\��Y�0�i����Y_,����f��0Ʊj�Pı�mTK��[tu�3J���n+5#��l�.v�4���J4E����i��	�&�Wa�0�6�fm��*dnhf�f։���!4vsD�v�t���N�Ɯ�&�	��;h1�ҕk�h;\3mQ��c�چ��J��+l��:�+2��d%��H|��z�ƃE@��e���7
�lbR�tV�6Ki�n��7k��I�z�[�Vi�B%�/��EҸֹ�0a��2�Fi�dۍ�(ZLH�W�.�f�)���8�m��Z�9u�nF�Z�tU!	q��4���a��W����l2����0��ͦ*����2��7J����c^8��RY��dd��RC��u�o�)���؄v�˯��_OC�B��i���3ZV^�2M r�%��[u[�VV�aQ�en����*9^�0��ۖbh��C#Lm]EW	+����6�u�v�H�f�AK4�7]y�ꝱ,.9�hm��X�!�m6Io.5ح@#���e�l )�ɶA+b��]-�uf&6�F�\�2�݃6mT���x��#�����)Ǚ����Fh4�����g[.��eғُ�����]���`Mم�Y��l��S�ub�1����pan�3`�b]���R�;��5[N��:��B�*
12�ڸ&׍��e�#F�K���45pQ��8bB�źl���iW1[��VP�d����ZM5n� e�م�Ɓ]sq�����iK��l�iW[jEq��դbg���DIj!�e"�7!�d��ibr����.
�qe���+Pa[Pu����g�*^q�v԰���3��Ʈn"�5��d-����}Ӥ�:w~���3u@?�?����CZ�)h�N�qt`�J!`�����l��wˑ6�,{��o�qc'�o�A5�T�˸�.t�}�9F9L����q��x�]����f7��8}�<���kiQ�sn��#�=MW���m=�vxgri,f�Ȍu���	�HݞZ�y�i�뤿z������}gtx�s������]�oU�m�O6�ùs�����ݹ��e�ȹ��СF�uڳjr뮨^��.�U��ֆ��d���Q�/��o'�j��$!���S�K�i�k��t���{�=�8�l4�ty�k�3J���NB�n]����^᪯n\95�[��]77�Wg�{��l�f)�i�<�bVe��Ln�e�rM�ǧh/`7���ϐ�<o\��:M�b�v���W@�K�gV��/[�=^jK4�۾ {ĩ���Ƹ~)�����m�<�	�go����ۛ	���EX;Îi\W�u��Ҙ(/ܷ7���V����9�d'o{K~�d�9M���O׎�!��Z�>��cÏfC{��TfnN<kU�ZC͍�o
fub�V� !���C��5S�4uy�gnY�{���	�RX�{	��_),�4M&Ě�e��lMN��Z��f���@��f�]�����!��w|�e7�:N��{E�=b�u�Y�rg������<[�4/u!�ug���/ӓ���s$hfʠ�:74Z�ܽ���u��F���[ڃ��E�bvY�D�.�(�v�`7a)���il�Q�N>͗��{��ٗ�XX���7ǻ8�[���eK��ߺYNj��zrsݏ^ �}nr�k����.�7Zsr��S�,�Y��U�Վ�����tc�E@����q��;�I�C��1N�����"&� ������g��{/ܱ�y^�=�-Z�Iޱ�؊N�Z�����\����"�K���(L섐1����ǏS��������v^S���Y0�xI��H���������;���ε�������u�J	�����F2z�`��)�4�;�����e����1g��d�4�m�.��ۤrS�T�;Ý�f�R+�Iv�({y��}��8N����l���=4��S]n����Qy��j�N��,D���=y��\NeeF�K�pc0�wC$<%��ɉ���q㼠�o�5o��]��޽�5�ԩ��Vpܾ��s��w���ӂ�{Ǫ�_��囒�1�V/4w���>ND�#E��;�
�GZO�^�^�Fن��,�Z;L3��O���M���^ ��+�;&���>~��WM�4+��`�5=�d��~]Ei�#3�T2m��Dy!�6�&XR��P���(�����9���n��Ł�t] žM����Cs�RQd���=�y��on�ӹA�s�+��r�$�8r��uū�w�r�s^v����ز���T�9��;}��]�wgW1j�����X�o����^�����Qz:�1�Ӭ[��ϯ�Ѿ���n.�_���wܫ��z�zhj{��W����{\��d��t�x�·�,ʹ�ه^n2�V*��3*�)�N]�D�.�u�a���x��xo[0VD��'�������ܗ)�w__/x	����q�<��F{��-��W	^�|������ü�nj�������M�Ҩ�N&MV�`*j�U嶂���M7���g�I<�编�x'��$�>�����A]=n$ӱT�8Y�پڬ�!T�	'�D��\;V�cF��C{��nc3�o=})L�z}�C�5��t�&M�������Y�֪78�#x��. p���*���l6t���i�^�������6�\�$i��N~<Ѩ���E�ӓ��帼%H�8j���6�G-�cõLV��'K�ub�I�0j�sCX����5���]H��U#�lY����[�{��$ àH�Q12&E�TfՇw0wSb��e��b� �T�K�t��x5��͇/Z{D���LSVd�,Ƭ:�h��J5�P7�M�Z�'��Bi�ұ���E_����cږ{�#�<�sݴ5Px��%���wޓ�3���3f��^��z��W�w���!̞2d�:�MV��b"��dM=�ך�@>/տ]��A����q�����q7�ٲ�Nu��lD*��0�]���/*�}���O<��T5��u��>Y�D��W�k�y�єvԺ^s�゙��^��^y>�����x{9a���Z^���n�p�No�������a�$P�ܕ����M�z2Xw��/e��A�Y�	� I��:��������}��h�@%R��^�h��bͲἬ�+C9w���r��O�ь�)� ��P�T��N�E㜇g�{̟xٳ��p��Lc�ZF���mEb�5�.�	�'J
ٻ3���D�{�t	�����݃`��LF�ly9��*8v�us�f�a�Y��#Z��w.�Ѷ���{!�a�F�����L#���4f�Ĥ�t���H"��ttn�15HV���Ӵ��e��n c�`��7xtV�'���A���<x�7D3�{"ɴm�B諗BC��1C��qj.ۑo�Pb���]֒�Nm�۫��\�P�ٯ7���/Ω�u�y���K��y���s��$8w;b�(�7�����oc�틎nm��6�N�@{�Q6��Rp�Dض7�rj�����=��px��<�:�Os�6�E��>�`m��)��o����sve��f,�޾��(�1�kն��N���'Ҭ�~��{��R^�����B�b9����n(����B��F8N�a�K�4�n��]�%�;��󻧎�g{%���i�`�7n�n��7R^E׶L ��@8���ଃ�Qb�-Y�A��S-���gV//YX�ئZ9��\�Skl�֢�Y��4wZ��I�S aƪ���vXV�3��NP��q�k��mT�� ���[��;᯴;�Ȯ�˽�;���G.B�j�||O�F��z���H�O/y��U}�����Y%�E�>��}��T	��[�/{�՝97;���~�}�E�M������{N�Rr���>�8��8�\�̦31n�V͢���b! �QSKa�­8n�ç���e�^y4ڑ�N{)!=˝y��3�iz��B��{-�����#�no?M��?g�"ޫ/^�>^��1.��v�@�2Ýs�g�P��fN�nhǇ��m^�j����Qb*nX[6f�t�"'e�ܛSBwNg�x�X�~�5X=��:KQu�;Brl�Ȅ��:�vo*�gD�u>��{5M�^����ɱ��I�Z�um˜ŀ{��vo�����C���ƍ�u��y rL@����[q�t�Ok�sF�>\�	}�;�̞ۈ��Ew9�`>�G�U�1�|�����8����ݬ�I��,�;��U�T�lP[.ÔM����9���/.N�S����ܼ�D�|��� ��4�v\����C���{ϗ,R懽;D�/��#]w�K�r�?f-��Z����=xr�9fc�UgN��D{�˶6�/�q�˜yl�Z����f�.m����-81>H��L�PX��gXuV�y츺 �7v���c�tL�l����m�%���s]f���Uޯ�l+O��6��Y�F""���Z�K,*�la�V�+��%~Ţ9��#̧�z:�!���R��88z�p���f����(��Mka�֌͜�P�ˤB����`�r*�V��Y8�WBqNa�݅g���E��� ���<�|sv�h�ٻ���Ӥ�z6�>����X7�W��هbywY�bj����c��ww��4�l�}��D�͂�㖖�n�dû�q�ʢ����Y8E��wTfL�;[2��n��[P���a{��:���4x���}:�vЬM�����"���w�2^rI���6[#˝�zL�Is\�ȧ���ҋO����"�p��m �[S"⩓���u�^��os^�d$(�Us�"rx�!7���{���ԗ�=�0~(���g`;i�:��3a�r��Yb�-?J<���k�*�n ^�'.�4f����uz9N' �ղ��÷�s�
��=���2�������Û�v`�v�7�{<r7��g�nI
{˛|���Uc����+%^C۱[���n�yU��|*�K��]� [t>O!�<�� �&<�{��Pa�Q��%��OJrRN$��}�i�b̩��Zs��vf�y���γ��T�/m���g���z	$��=���zPb����E@��+ݪ�y�;���w�o��q�г�Rm(l����x�2����d�r
pZ},��p��!go��]5z]���2LM�ֻ��a^*zw/w��pk�2!����
�zl�62F�1p*��ٹm`�A�
���'}ŎⅢw^����D۔Y2-7�Æʙ�"$w��j�!w�s�ŭ���6a�s��y]��5�.�ش�Jp���'$FjdK�aD-��6�*�-�;��ם��K��̅$Ǵ�����78���/�	��S�wr��6�એbcu�q"����.0��p�wb]��z��z�gW��Ǔj�zy��z�`IU��=��(�7�۪zg��<�	j4W`��zyk�5w+��L��h���(^m�Y<��ٞo���)����piP����e�Oh�l���W{�r�gg�~y��-ԙU�|p�����([*�#W���F�M%ףSˀ�}�ͩ���z����Kݝ�T��D�� ��S9�7�0�,�~��*{�e���nv.��v���`ڰuֻ���.��7�;=6a���z^�}N�A����N���9�e��u��]�`;fP�h���{�O����(��i�gk]B��vE�ՠ�/�9ᚸ����c1���A��N5��C��"�����c+KR��9��F��wO��ɛ��篰x6<��Z�a�W"�h%����g;���|{F�aXbS��ž�sC�9{��|�f����\13� �=/g� �,DD���q{���2>l��y\�i����7��������L����9��*��q� w{��[���%��UՂꉈ�D Կ"���!.��b��/{.�V���-�S�&�%�De�n����X���Ni[/1���T��&f&��z���}����kQ�7sC%j���˲�V�C�Q�oqd�n!��O������t��+�L����;ػ򂾓�s����ۋ��:[Ź���CG��14+A;�	}ώJ���
�'�i����e[oL���#����F����1>�7ꪩ��8V����ꞳС���/y�T�����nW�sd�	;��q�$!�ߕ���<���k������J+�uّd|���}��&,|s�O�k��g���챞ɺ�}9��#�;�7��#�w�Ҫ��v0o=s���M3�#em��2���&x��ٱ����`�6��d��t[1����aXGrk�!Z�"sr��T�Ǒ���.�pq�ӻ���'�@�+�ٳ�k��7_Q���}^ �x*=��9�����X��#�'��M啂���5!L�uWqZ%X�Z���;�#�<�/���E����f�Z�u�w���$V���9����,J}��I�&nol�*6\ẻ�5 �� �vCfo�Ǖ�;�RXL���z�='��%w,}3��p�B�m�g���jQI���혦%���eo��:��/���-�g�����򛏘e� �iz��F�?~[�u!�y��%g�;��?'ǲM]�ݯ9����w�����X�G{�X�����i5�U�K	'��9��t�Zi���fT�ݰ���r�v6Jډ���D��l9��l⁢\��ZiVF�eӝ�Fލ�{����3o���]Y4��~<��᯹��ە���m*��4jݥn+l��0���$��9l<}�L�B��g]e�~��5��<���$A�W�=���' �>�����<�<j{����=֟w�sɵ{�X��~aeL�{ �X���<�v��l]��p�����0�������hQ�-NM%�+�6���;�<����ًFp��';�����<\������4�H�F~�3���%�8�Zs	a�ϦN�%�.aU@ۇ0%��θ���Xn��_�L��d�4���w���41�����Fx,�=K������΋	~\ν��8Ap��Z�Ά	�S;���msܧ9�{�_x*s�x�HŜ��M������賃����N�7.���GW��s�,T�5���j�F�U�ܓ� ��i�3�ْn��yR{,�Q=�,������o�:�nj[p�����=�ە�Ѿo��
�����D%�^��Qq��=y��nN�ݦ����up�l�Њ0�3
$��_0*l�<Az�-Ѐ���6�2k������������Z�ҕ=��4���*K}�0-�{z��{`w�v�T��m��h����i~^����$ON>��H��@����x>�	��x�����Z��/r�"���׏rہ��霴F��^Ĺ�����^�4��<��1Z�Ѓ6�:��������O��
	���}ƿL8jӺ=Z����ݝ^H�w�g��}�۞.x�o7z.X���̔�úY�T�3����=K~��<�^j��(b}�8�}vgS��@�p{,>�z�s�e���
�5Ö13TS�p0�9s["�!k/v.����t�[�s�4N����� rs�`e��u0���^�J�K�g������`#���t��Sy��fR�c5�'d-��{�Or��v�:n��'��ߌa�<R�lh�{Gf��5��3a�!�\v�W�,Z��w�3���#o �t�Ǧ�� �V�n�ч� PMo����=�U	y��e<1ŕ�Ea����`��Vh��9)An��������z�D�Б;r9��O�Ӫ��p�{��~��09���;���t�t�_d��
 ��/���=��Y�gZ3��V�� �.�Miu��3Mb���mt�(��j"r�8U��#*\f���M�op5�P�3�b�Wq�.j��smT]�ԅ�mkt�U3V�)��1��.[��I�t�Dp��6)�;M�9��t�s,�L7s7S#���p�ajRZ9K��s�]�@�cQ�k%�W
��4��U���[ saU���]	��V�%�4P��w�K��d^V]��l%�̖X1-�I��sQ�WZ�Yk��)P��)53,ns�Z6B^\0�3Bֵ`�k��4 ɫ�ȇ4�-�қG�"8�5�J7@ckp;Esx{5�]�,�p-u��1Yt.&�a���5i*A�ԗA���8c���B[�l,�9MIK�A.���a���6-(k5�l�P�X�,��u�fQ��R�H�ՌBh^HuҼդ��)��4�M�Lb�4�
Zʰ!���]�&+e�0��k70�8J��u�v�x�!M
��
a)�&�J�4[�96��b7�]��5�u�F��+�	�43�mG�#��xKf1f�!K�X���Z5i��Z��H��:����!ZJ"���a�"�:���4tLD�cr��Wj�h�k���\-�c�7f[g^DV �T`me̱�jV�v�R���.R:6�Ԋ���uXZ��1-,n)fx1&f�ڗb�����&U��Z��K-����lR�����rI�D�����Dh�X��0X��5n	�QZF�l��U�`�!�Lg��Y�X�id(�B�eV��xF-.�X씥&�.F2�������5��#-��1��r�6���[-auK�c�K`i�rd/��Zd�����Z�!��XT�^	A����S�B���h8���mFj�54f�X�ct�L�f�x��j���K�M�t5�@K�bi��n�4TpԔ��l	W2ض��K�H���ƶlk�TM��h䔆���h���"J,��]T*: �0ŕ�U���&�2�`��cJK��%P]n�	EX�+��g"���{�=����w���_]8����)x�ͻz��1�g�S�I�M;��37H\3s�n	)��"L�oy,�{��B�Y��F�A�	q�/a��Z:�"&�m��L�_�<�O�n˼j�/�P�<#�o���>�;�<�yb����Z#�t����E^�D�[��̋�w>rz� ���-A��i��h�A6�G{穀���|��7�E>м��q�+��I����{n�i�NH���/h�t��n�+4�3p�ӃJ����ԧ%;��=T����e���nSQ�$���i�:w��-�)�q�cܢ�Э#(;�^n���j4��9c@C�Ԡ��w'���.A�����$�*=�"��a����kK���[�9��ז�̚$�H�[���eE��#ۻ�A�t`*�ћ�J�����/yO9�D�1���=��k����d����o�[V�1�r٭�9xf�P�ϸ����y'���j�F9M���Ԓ�%D��"i�<��f�5�K{���~�hY6�4��fy�_���d�p���1R��>w���FGx	���d]qo��ۄ��G}��s����;��r���%��N?m#[���bs^���u�t�\�������f�5�w[���knAVlܕJːr~���ޞ�&/Y��W������%�����]����R�V���Bv��'c��$����ELܶ���8����b��8��+-8�����f�l�U�T�R6d:hZ��U`{̠�ڈP	�]��4��؍,Z���X�]
`՚�M��刼�5�õx�������bR�b9�EV�3��X�sqK
�GMR*ʕpV��I�n\��F:����6�[EA�ڙu�X�H�N;\Z�q)n�%m��Q�۵�0��L��aĦGL�C���ź<�fW��f&m�1v�4�%���5�@�"�ү���U�%�*oR2Ҡ�6�_�^c���Vvz9����OJǼmO�J��c�7�Wc<1Z|��2��?���d��{�}E)@�1e���JX������%!PBXRY�9���������بY�䴋�Eڛ	z���fC%� l>,�S��zi0^/f0��"fG���� �!�
�̌�V���N�0���>f�Χf���Yp�}����I�<;=�����b�q�X��	�%��K� �º��l5&�e��f�D��Lw
�,�µ8f=S)G�̩X5�'d�)��U�/�q[+
�]�=5����'7ř�xXQ���t�K�ħ�	�DIM���� V-fgt�wg�Q&N�+�.�aG�v{�o@�i��2�$��B��̀e+f�(�%�mЀ�h����f�5��k��;D�Wl���<����;9����YB����L%�N �`���̚$�sK���Wc/aS�	���%򘑽�K��#ZH{����}{��/m�����o�)��I��z ��Tc�\E��i*�k
}���li��>UhMϲ�=��'`��>�SS����Ǻ��xܧ�{��"q&N���$x�����(sx9�x��\��xC|%C'��=�d/���l(Zl�k��G G���<�a��}��) y�a&�W�M%�L̊��Md$�f���+FI��
Ƴ��E��a\�X�YׇG�М�ג���������#Q��(XIf�!%�o������:<'g�?�ҋ�c �������U�ş�+��T�	����P��Y��V���D�bAf����g���t!3k�Ճ��e\V-Fb5�����gr@��2^��v���zNϬƮ��2t���+�t�-��\<G��,wg�X*0��
�
�!�$��O��3����@Y�$��wd��,$�e{`�4����VjfX�<,��!ݡa(�(Q	L�yE��.%�#O���ZEw�^�*�^�ٮ��(x��2�&����l�5�}�I�O&�a\Y��"j�\�G����e>���Z��şh�c��5��8Zs��ń]ӈ�6�%;z�e UN��=����qK^uW9���������}� ͙խo���0�$��͙"ϰ�٦`�Y�>�
�HR�Q>e
�3�����h�5e���K<,����K51#0Q;�.a�lu{�&��3#���D�V
�(SyO*ƳƳ4�5	�ǳJ����}�Ka�G¯a1��Ny��-����1+6k��R�v�E���0[�k�FY��;�(B4]�i�}Y�=ZA���-,	����2���~#�A{*`c\��֤2�& M���}�(���\�1J�kI�l�'�*.�%��He"_!/����{b���͘��df�ȯp �#e�Ek]2�k�3n�j����o;�~"~:�(�cj@����a�g4�<`�63��O�3��;�u�)�\�ag_��53�fAFk��	0�\V��9b�[�����>'��qN�ḱ��wL��X�z�`%�̈ Y\�ѽ3�I@�>�ढ���b)�	L��<D)�>)�=���$ydEva�*�a�Q��M��m�����w�@����e�W7SR��fӺ�޽�T<,�1�������f4�櫝����$D6�i��g��C���!�8�*��ay��YB�ʧE�bb!�"��i����<l;6k�����65��C]�c �\����r!։ހ�tM����ΏI&t�+3'�V*,�a��0̖g�U¸�dY�J�S1D)���Ed�
�
�S!��j3_~�XI�ms��:En�x }����1�5�Fڣ��5w^�����ړß�Qx��5�|2�'zvV�,<y��ׯ	�Ώ�<��Ɖp)ꩧ���'fo�y_lSQ��}�D�B��2}b��d�f�e�>|�׆��Ď����S����<�v�����K�@�c��`�4����VIe
o+"��"�'��*��Ko*��.dM�\�h 0�6�뮡�)�@�v�M�H�ڟYG��Z����pg�q��$�nG�/d�7[+˒ab]��F��\;/���2�M*�m����`HP�lcc���9oĈ�L6b�n2��@��\]ʙR1[n�����h�n�斍�͆�Qـv��
�M��a��\CF�u��i(B7CAtRg����1N��XT3�9KaC��Szk������RQLUΎ.��a�B���R�`Xa�49������Ü�$������Eȝ?]�ȳ��{O)H[�;����|�ozZ2�̔f���<��)��\�7��^�S�)��P��T��Sg@X*C#@�,`�SYt5���R��k��^�#���-��!�1?/�ܭ��TY��}2+�F^*�CxfXQ��+j[JoQJR�$'�ff��>��k>����3x^0�n����I�nHYB��3)���d�eb^0�?ʝք"f����x_�����Vx�|^O���S���a�vU�+I���d�P�����k���6[�:?�N@����~�aB�h˝��Qg��TȰk5�gd��;�f��Ȣ�{�$�L�"&ʉ��
�.����xo�0�Ik�k�<,ܯ����E�e
�ԕﵼ�Z�Pq���%v3,�	+��2�݈��A��#��%�L{��p�7�]t,P���1Z)0�M�P�k<,��EY%��g�[Y�� d�xX|di聆P4���/ �e$�-�[k81�6w��~Ȏtw@V�u���un='ރx��e�F��������d�x�BL�$�2��<u
�g�}�:@̤�n�U��"���S���Ru��nE��,��T�UtTM��Gv�F	�tP	��g��-��i݅ji�����̑e����@�h����Ag��G�՚�pG9��}o�{�ks�5\޽;<'g譖��eW���V�N�I�'_5:�~��~��1����d<$�nYB�ff[��Eh�7h�cY�\�dՔY�±�02߽-��
.=��p���	��"����$��d�l Pgӿ=5/f��e
Ƌ���|k0#}�x�痗��ˉB�6��!�L��;1p�R�t��[�]Y@x�<-��5���MRR�'�<:%����(�P�3Ұ�Y%�禵$P�x��J|f4FG�Q��
<��3�)>��r�f%�`ۻ?Eh�6qB����Uf�x``M�����Yp��12^z$�����S�*����+$ֱ�M�)Q%��m �7"��ܑD��Q��z���T�Fr��<(�	)\����ӻX(��K�d�����I9�DWL3�%�-�l�o1�	Y����:���i�ϧ��Ԯx�M�	��qn��+C��5�Ï�Q�,���+�p�:�̖@�o����0�yq31V*/S:IYS� �l<-��������}-e
�xh6^Od�"�����YS��L��\y�N���ו�SQb�I�P��5>l����c��kE�IyO���ry:�y�Jݳ�˄�Y���
7G:�imi���-�mV+�u��"g^�͸�7H�IR ��)�,�.�8�h�6v�5�����k$A�Ca�
W��MG���y��-J���f���~9�x���Y!P�Tab�n�_���YⰢ��^O�Y�}n��X|}��r�E/̴(rff�^����(Y��g5�	�P��!���r}5���#����
�Mb��?��9y�O�)o�3%��z�|���9�i}�D�Ƌ���$�����0A r\�'r<Y$⊚�i������	��Ǣ��}�G`�>�Q��a7��-�5�X��2���o=�N\|��mW�q�K��=�f]f����'�������>qF�s�)���8��٭�$x�%�4�fȑ[�2�"$��3*�E�»����bԐ��`i�ڊ�Q���ơX�xQ�g�Ʀ��9��$�Ȁ��7�M���&]��lr�M�(b�[@H�''?�:l%�N��Z-s�ztM$��zj��d�b�YB�2�z�Ν���E��d�>8w�V"�R"b�35���,���z��q|2q��V��L���k(Vx|+0��
@�@�G�Zz,���Ѫi���ؾ��=5/
�*&�5���@ӛ;�����i��#�U	D0����A"b^��f�#��ߥaB�O�����y ���d6	��}��i��I�M���ݳ���O�?y����t~(Ԑ�}���P�x[3�U�X�M�KXc8h���� pt���t"�����!h���r���n!�#-x+Ww+�J|��$� {i
�,����6a+o�{�JM��n�B��
P�M�`�����a� ���[�T���v��ֹlx)5r��1Z��&��s���9�n��j�63\t3�kŲ�E���#�u��ڜB�8Ȑ�ԍY�p:�Y���II`�C;�H���S�ܐP�\Q��Y�1����J���ut�+M�v�ݍ������C�,�sW(�ŋ��0٥`i����:�5��cZ�pR.� ��L{�����7��Q1swY�;$K=� ,�T��N��f��+ӗ`p�Xу
$������.7��%�!��q���+K�WF�l��3qb��J8ۘ�5cf�Ƅ[`�s[����#�n��]g�+UV[3$IHL�Y}'Z�0���YZ�zN��w��!�+�
�ͨ�|^�w�G<3ƻl�~9�I���:��K��M�#~�҅��~�M`�7�x�Y��r�	���������[p\�t�1%3�)�w�Ec]�zk�d������(Y�6GO;U�N�g�ЖHI����"Z��d��ƲV��+I�;�Y�<�xSAf���xQ��}1<9��^�T��tٖ�u�������d��H�^��V�0^2+g�h�4sm�S"Ϭ��u�ЦB�D�xbm���]ITYf��m��fj���,M�b9�s�4�����RӪ%��-,���b�3�)2/$,�X�q���a�|/��Αu�0��#�b�(�D!LkL"�wS�=�bL�1&�;(�#�����Q�T�{)Y�b}g�����n��}�$��p�	M�1�b�tI+��$�X|8�r�{viyTK�ˆ)�FM�M9��K_g��Ur4���M����h8��~��e^�[U��%�]��xTNi8�ߨ��g
����>������S��{�$��"xN�퇓\_@n����^�8�`ѝ���χ��cs2I,(W3�V�0_��P��!��2�D�)���Y��I�4�����P�/ة��H�y!d
�L2g̍�kI���G��ۭjQnRxs��,]��X���̖�ޖ�E����V/���������ڂ�J	)�D����m�n4Κ�{a҂�InT2�%���n�bp��wV�3#��'�觞{v+��z�Ag��X�Ra6����nV��(�x��@h)bS��LC��YDi�9-�g�Y���!�6F�oM4*�w�Y�f�`��ꘈ�xP�)�"&kEFM�T:�����*�=��dnuj�쭭��ġ��T��Vc��1�"Ucs�U>|�d�&�Ol,��}c�����N&����y��.j�+E޸�o�]I��4�5��sZ�P���܅H;���{�����蜌����V���sR�GU"�����ۊ��^-{�����2�'n�I雍�g-�uߤ�O�Q� ��3�#q�l�/�����|�x����Y�6i��kN�;5S.cn3��	nl##.%�ǻ�׳Of��5F�Ts�'_���}��M�8m:�?�z�0*�ն���U
��dgt�쉱�*]�v#�]˷�ji��/@���1[z&�)u�S�K-s���;��r�Z:nYv�9��Ԭ�����Mh�<T����z��b�j�{k�o��J�x�h;b�}!���O.��n8��i۶!�Q,�RQϝ_,��᷵DA�u���Cy�:o�嫚v{r����mD��dGq�^���7�*Y�p�/��ez/#�p��+�S1�ȹ4�T��v����9��wBOa�.��u�1D	38+��\�j�m����eek�ww8��ڙÛ�ێ����к��e��t{����׺�$e������g�@�V\�<�K�=Wi��O=��eqp@�� �b��U/��7�e�}f����թ#1���Y�oON��ؽi����}�2�J�^Q�Yz���=�w5<0�оO�Ut�N��#�t���B4���!in��q�7������S�2aV��Em%�6b+N�z��%�f$S��o���[aS[9�͝��b�1Q�DS�g�2�~���{j��h��g2U�q^� }�Nm=,gn"A���͡������F;���������C�<��q��{�r�:%GGj�]O�g��V�!F��(�MN&�۫�0�L�s�j�;��]�
e�����N�=���1�V]�RAgI1���}�+Xjd�/a��ꃷ�V9��I�s��qW��v�{��á{0�Iǡ�v`�T��n�u�>�N�v���xe n�9v���"0\-��ǧN�g�Mˡ[����x��7�}�	;y��ţv���e�}���)˼@)�0�:ITĩ�y&�������t������˩��)	Fo�������J0�m`�w���=E٬a�Ym'Q����a�V��]kݡF�q�_�צ���x%^7���듞�+R��4��n�h�&�1�T���k^K��rRoӲL5�b�?W���-�0������ޘ��6���M�αd�Qw�3�P�/*1/w�,�uy]����Ǉ��{W'�J7���/�ft���0�i)g�v��~;��W�'�����:Թo`�F�ŕ~h�%蔤IQ1٬FZ*��0N����([̒Qv.��ѥ�X�L�Λ��=������4e>Dk�k=.��Ԩޱ�9����n����wΡ��~�7��N2�>�֞�	a�ڠp����΢�6�u*�Xq<f�4a۽5��M��˞�!��:k*�K{4����N{�*]+p�g$HU\�|E�#�w\����8�0��{��_�T���(�T�;ֻ��R'����T���/�����<��))Cs���?66eq0�3��Wޯ�Kg���Mɒ�!М��
��Z5�7��7%(R�9(s0J7
d�=�}i5rry��{�R����o�;�}��@9'�d�I�J�9	����ZD���))yx��<���x�m/����ӽ��rrL�w9	�b�@d����J_g$]�	B�d���� ���y�p�قQ�S$��܉��s�����d��2_g$]�	G;߼4)�)(G��Os(�I���.����鬻�;��9�l�'SB��i����Q"�ڛm�ieyn�}�-�s<�m��m�}N�y��={�/I���!�����}֝�s0��d��/��S�׼�Д!����=���b���4�BS ~�%܉���D�����Z���)��(�)�y&@t>k�iH(JDJ����U
����{��<��(R�S�/�׼�Д{�t�t!I�L�99	�`s��Zp�%.�$Nf	F����}֓P'!7��G� RR�׾�4�@�`���=a'@��rL�=���9ff��.���:�-�}뮴%������Bk0B�}��;����K���`�y"d��^h�R����>�: ��'��K��o�N�f	F�L���79	�}�.��G� �&K���`�k�}�f]]u�WqtZW5�z�@nJJ�r���5Ҕ�!G�(k�}v����GY�R��2J������`�n�=�%�#�����"Q���!�q�L����R!���Y�>�W�x�	�꺳P�<�6���G��jsR�,v��>�F����"�C��).�"bd�1_�᰼�Rl�����O��(g��L�G�ӭ��m��g',ڑY	�@��xJC������7'�2D�r��
<��=�d~J��r��I�{��ow������Q�!�y&@�~�y�N�9��G� ��r!���S����%5
�Gp�s_��
w ��5#��{��{(��T8�Fds(��:�mѷ���K�FV�V6m�ʕX�*R�"$��.k�;�I=�1m-�[�����;�=�,��`��d��2_'!����	G!��g!7�!G���;��=�%�rD�0J<�rOy�����0L���f*Q���L��y��;�9�%���M�Bw����]�܆��������l���
��%�G!<�T��w�:���2H�R��
]NB���!rO{��i�_�!7��G�*R����;�9�%��=� OӐ���o��	G 2~\z��B�������,Р串H��I"��RK�-$�!9�	F�2�}k�'R�r�`���I�.K���pӹ��Q�!�#�����Os|��B�}�nP�y9
y�%~߿Z�% jr��J7�_����#V��=:{Ǻk��x�:k0J=����:D�)5�}�w	�b���^I��9
u�o�	Br!)_g!5��G�o�Zp<�%�!=�C��?TSЅ�s��֐)y9(o0J9"d�9)�}ߒ�M�U��rK�z�s�ry�	F�2D��rT�s�gZ�J䚓 g!7����k�|h��NH��B9';��v��=���b��d)K߾�i�	��)]�d�ɐ���O�'����g�j|H��7�G��]�@>�\�k�&N��s@A���#7d��}��<`Y�b�L�� i���)��E)]�r3g-6��!m�,
z� &�ܩ�.�f6��8��B,�P���vG\56m͉.�B�t%V�Y��l-V�f	mHQ���+�Z�5����LRh�\��CkG��ɯT��<���ƨ������i��[d.�U�eV��V��8ڎ�ɘ�bV$�:6d^�k��W�˭�!�
!�!� N2l�L��s(�o������ef�E��,���=�_q��[Ș����Kx���Z/�_>T��[�=sv>��y���:��$�(H M��ն�M�f��F�kj"��k/k*f3p�횋\2��N��o;�{Mٟ��)���BQ�C$���������8h�����C��(��=�Z�i(C��M�Q�I�K���pӹ?�焭�'�`�u d�����Ns���Z���ܙ/.RrO�g N��ށ���:�:��)(]NB{��F�2P����&����B���Cy�P=@d��K��ϳN���PI�2_�9	��w��B�r$�i}��w�%��iCr{&C�r�79	�`%�d��ψ�}�gVwthLֻդ����`�r�7&J��<�����n 
J_'!N{�<�BR��d��/��NBy�	G��ύ������b���9߿u���r�d�	��IN@�	#���hk}[l��I�u޻ӸNf(��I�|@{��GH����y�y�}�J<��))^NBk0R���ܴ�}�%�rP�0J7(d��\Ѥ�NBo0B�`2>H�G�:�����Ӹ��(N�2JJA��}�s�/�c5�W��u�Ӻ��<99)���E�!<�������ܔK����(ܟA�����}�MH?NBk1� 2JB���֝Ȝ�����2@��';�5Z������rQ�`�|'z����õ�6���:�S,K��vE�
b�s�X�h�������]�	Vh_�'��u�7'$�CS������:��h�R�9�`���&�2]~�<���`�nD�))|��N��|-���.���I�%���`�}��� nJJP�p���9��Jry���vn:V;�ɺﾻMK���`�{(d���~���Y���G�W8����'~ǁ��k�q%�غ�K���:�P7�*��=��6��I��f�:3 �>+���CV�ی8�ߌ��n>L�؋��S/�NwI3�}��L�1r�яl�Gg%`�����qG;�5 Q���/'$K��s��%/�����rY��~�9�7+�/�	�`��2Owֹ������;��?f	G#����䤓�~�llf#�z䛦��N�=�D����)|��=����	G�9&����M�*Q�~����))w9���4t/3��)�u��٤�@��&�h������Ϲ�w s0J�.OJs�~9I�����e
�5i�$�uގ�%�rJJ_c�:��
y��k�����.K��!��(�W$�߼Ѥ�NNBk0R�`2MB俷�yi�	��(�P�)(>C�NBk�w�iZ>��T�9��s�[9t�>��R�G:N��u�7%%!��'���n }��u�j^N@���$��s���\�_u�p�قQ�)�rL���Bk�}����d�-/�����Q���ZSr{&B�9	��;$���Oz���3`��U��� ���5�k�R�,�T��f	�Z[���%R�C,e��޾�ow���'��Q�$�L��_}i�'3(�%))|��=�y�}�J��rd���&�(��y�h�2�IK�	��
?@d�g9�h�y9
k0J9 d���{�o���M�Ϻ����Ο�ӥ�Y!z}�������V���|B`�%% rry�s}�zp�$�u9 s0J?@�'^��% {9	��J=��I���7�N�f	_aԥП�:����9	�Y~�Z=�=��oSӥ�����סW�	�b��߼�@nJ�S����Q�I��]��}���`��ҵ�m_;CX�7�Q>��z��𯔟�"g!�:׆!�#��`�j4�����V7�})P91���ݐ!�{�{�X��P)3P��=4H�#���˱�b����}Vs�+[�u���&�K�,�w<�=�-.�p�J}����S����������z=�ܙ�X�q�2�����;�<���L��� ~���]s�iB�`2����]圁<������ �h޹κ^�RN�NI�������N�� 2z��4��NH��% 2O r_���Ɲ�� ������=���=��7#��9/�g ����%��ߺһ�����'3��I��v��yq�14�UOL�/�����erJJ@�}�i�'3�P)�/���_z ��߷����II@���b�u�}�Zr'�d���'��y�u�sF����!�`�{�nL�Ϲ9���~���'�,������K����v�V:�[!F���`��ɷԓ^ϯ��/$��%SSJ��e���I8� )|��;��|f���Iܙ+��'���{�{���)){��=��$���λMO��J�9	��
;��JJ_uϷ�w}�%�'$�C�䦾����;ã��g]���BQ�IIK�By��G���rr~N��Bd�� f	GrI�5��% }9	��h�I�K����4��`�y d�����'��<�G�?)�:�O��)9#l�	���}���ŝ�w��ֵրܔ���NfQ�Ju�_s�'r�9w�%�IJ��]���0J;��:w	��rL���	���iB� 2J�����ﵾu�����NO-��'d���_��Kw;L�z\�k4���J��%��t&	I�2�>���p�f(Q�J�R�9��{��`2N��g!<����u�7)IK�&B{��7����23������uoB�zWu>*��&�[^��9>���y�V�VB����q�+���%����ѥ9-�W����O,c<�qՋ���W���/yhy	^��;�C�rN��ɽ8Rǳ�+"�C@��{z��A#��x�$�z��]��y9w�%�rJ`s����, �)a:�*���d���
;��=��NH�u��BQ�&IIH�9	�b|��h�k�@n�2_'$f	F�rMw�ZJW���f(Q�Hy&K��˝����(�2JJG��O��?S�"Z��d����D�L�- h�9��ݴ�c���D&̷Z�Z2~9�Z����������}�J9�nL���&� (�}�ZrR4����0J<��.����ԯ����V�`2JV�;��f���b�f	F�rNI�?�!>�j�!G�IKÔ���g O��{�:�)���^���=�!|���0��d��-%/'/��13�y�n%��}�i��`�y�RR�����<�G�&�2_g!�	G���w�w%%×X�NB~N�������~�L�	]�����5/Ӑ�y�Q�IIB���֝�s1��2_d�NB�����%!�II_!�K������G_k�p<�%�C!9����5������5�%��]��?�?��Ѷ�i��x�|���y�Q��]��rP�s����(��nL���&����}�Zp����=��%���y�M@�9	��h�#��:�F��9Ͽu�p�قP��9&B��Yҳ����f�f�4�����o�K��))}�!5�!G9���=��{���1o/��n��}���24�3��sדk����M����4^�1�C�
�C�v�ّG�ng�3���>vF������8L�����2��T�Ί']��i{����3���|���E,��a��BĄ���v���q��V��qv�M�.�E�6]�-�Kak�R���,��:i-�ڄPf��:�3S@i�ަ���b�f��s��λb�(��u�Ŵ�����0��^��lٛB����.-,��a�M�kl�ʶ֩��T�,�� �-�]��ZĎ�TM�+\�F�.�G[(V�PCe��"h�QRb��{0(Q�e(Y��d\O�JjFu�����2�0^�����5u��Cw�n(��9��[�`��rѱ�,/ 8��Y@L���T� �s3k7Si��rd��`��m�C��׸��J)(���J����W��&`x�@k�f�)<�^2��*�hLy3�<֣�r(|B�Ĺ`�î����7��� ���JP$) ���q�-�O��+K�i��lÎ���s*���C6��b���+����;1�3_ʰ��d�Jo�D3;VN�:	R�0�	`TLҿ� �,+��ՊGX^>�2kvk͏'3#D���Q�9��T=� �^�[_|+<9=k�A�\�AB:�2׸׮�������s��H��z)y��ٵס'�Ή���Bc�/���r ��� a�y��D_���1�~]&b$�DD���7�=)� �^wS�q�Z	����>�Uw��X��x/Rw/�b�f��L�hk�~���/>���K��@��d�+SZ�-�ZY�MD�XhGgf�`L\�\�����A��t�.��_�zϧq��N^Lw|��x�@5� =�jExr�����n�rHf��+Z�C3�� ���#��{���>y��qtMG�gu�������»�r﨣2���\B�Ul�}7y1�
1��-��&]Ht�0S�eJ��lآ���fs~��a����v�i8t��V��yM��m.�cS7p�&}�#��>�ih���{>��H��dTPP`T `{��\`x��ɫQ@r	���1��By�ׯk�L&hJ�HJ�F���u!DL�~QT�}~^��_p���%������jZ�9�)F�dq|��\� ��K��&,W��`B���t�3#��#���Q��y��a5I;k��3��������U��L ���Qݒ���c{|�N���������;�]7�~�~���Rn��6�����O���&����|���_�
D�������a��x޿��H� ��X�q^��އ��e�x&]S��p��0�&KVnՎ��Z�����e�M+�F|�ξo��*���
m(x�q�&��Ems��3;	cჳ�¬Xa�q�ݗ>� @}�<P����|+=�/b򤌑�/�H)D)����`;���VW��}��� ������O�WLּ���'':+��>���z`�s&(��:���w�&0A/O̦j�}�ɩ�b�hz텇� ���M��Ձ�g�刈����$��ڕeo��xQ"Lx>� q�֧�׉��UB%q|Z�y���i��5^���g�4VVH���@Wᒸ��Y��tEu�75���]n��*�Q[�G�� b;C�l-F${9l[����!R���T4���!�y���.���ɔ�M�E{)3 ��]�DD�"$Q�=K֞eN��u0&���q�$^����������g��_,��&a��	�����$p�ζ�.x�A�,��EW�C)�ߧ��Y�?^��h�e����������@B|f��`�9;�^Z�җ�ߙ.���:\),�3j`tj��x8��\�m�Zb�)d��y���ו�4���Ǯ�n���&^���"�{���z�����EtqZ9�F�{�f��!p���hV��3��~3N.ў��H��A�K729*<�a��3^���-Z�Ӵ:tV�z+�ΪKd�ϑ�t��¸����搜��~��	7s���GlU��\���!�,+���Q|s�
�"��u�A�'3/8&�Z�A�o|���!OlئT��yHd���J* �&�����>E�'V3S#e]}@��D����G�u���6Y�˗�jf ��JIr��wOc�P*{@e���ӳu�'���/��}Q����$��$��x�@��%اs�z��fț�ӿn�a��!�|ʒ��=f����_C�����ݹ�:���)^��p�)T���x�7ڻ���8�@�o
���}�Q��k=�,^X�����̙0A�~Tԡ��E�3���M�C>�L�P=��O�M�!x�w�~h\ �CP��Y���x^Y�8>{��n+��+1YnڇZ��0��;F+�m�ˣ�٤��)���s��l��ROH)�U4�������WSiv�k ��8U��d �H��J��x��}����t}�E�T�I.���ݕ����4�}��}8rs���k��P.̵�Y][5���O��Y]�`�� �#Z��tyqa�w�f&D̩��)�6�!�{������ �f�5��V$�]d<ms�k�ҁ}ՑW�/Zf-A�:=1
`J�"��gl�ΙC:3��W|����|�G
��}���5宦�3"���Ϧ�2x����b�Q2�#B3�35J�v��"�,����}�A��.u0�K����F��S��ݏ�_%3	��w�.6�l�R&��^f2��Wa�!�S�˂��S%`��y��F�����*5��M>]��؜I�ƕ����ttp�i�l�1���	��G���ܘ��F{_��.NEL�{�&���]n�n��͏��ۃۺ�-�_��}ǈyu��ƌ���#�Yj �m�d�v��?��&�z{�����֋�20S�7B�N�t�m��M_n�T�2�m�kl�m8˾�7����7�ٙu3����s�A7xqf���O�x��jA��]�Li�X��5w1�ˣ�uڳ.8�̑��VpNy�2*刼����D̥�dY��N��3yZ;�+q�ݳ��Ρ.�_��o��ed���s[Gf[ι�
�rJT>ͪ�[�^��{�|��?Q3�w~��s�P��엕2�\��u�U:�nb�"A�#�;����LF%Zz��a²�oP��B�/�7�q�#�$v=���ȅ�H�ϽS�G�E���m��\��'��1�NdD���u�TSt��ja�{�j�6�FM�d�jw؜s=�*u����_�,m6߬�]I;ki��{V��ۛ�ݬqSp���V���Qw�Y�SЎ�"���+&�(��C�Vv^��f��*3�.��'�9��'��n����0Wk���ޛwӦv�5FWD�ɒ蜾�Fo'�9^�3�2��xyW�/u�v35�Q̊�U����A�%��זIH��
��)�DwU=�b�Te������l??b�t���+�B��<EtC̺��O~S/I�qf�/U�{&5�S��@��-�F����}�E'��t@4py��g�x���(����-P�d�re���s�-�KVD�7wJ$R���ؓ�P�t�v�r0�S��LI�*��h�$��θ|�n�������2�Uilrk�D���]��p�qe
�s%ģ/����1�I�b����ڲ��6�P�bXK�����@�jP��J\��L.+�oPeqk��-֔Y�PyaV:T�٥�6Z�c#cvm*J�+R�$�Z�Yb㔔З�-���Ĩ�%YNu�iF�b�k&+
VѮ���.fVe�Ҹ��bu(�f���Y�4�u�Q�T�p���Mȗ��M.	DfWR�B���لM�106��˭h�.,L��$Β��(��0FZڼkvq6�:�7*�;Y�E�fT¡H�H�a�BƄ�C	)]Ž����5�� Tԕ�MV�J͂]G��p+r��h��)H�\f�����i�6�%5���J�!mYpR5CZ��R�n�VZ'4�`��#�ց1���*�]�s͜<R��	�&u�`ՎִJ �,)�Q�Yt3tB,��q�C��Zق/⒦ɨ��q����a�tX����-�fitJj:���4�k���8�+T�V�BR�9�үY����:��9�i��ciJK3n �Df�F9�#@�	�Zi�k��k1fy�\eh��t�#�Qf�)����g8av%V�ku���r»����30�v�Mb2�KR�T�+58�X5Fe8[�R���D6�ݻl`!5�Ļew�V�FLSq�5N-5�w.��K�P�f�B��z�X�� e��y�Lذw
&�E�@�����&��%�1��%�L��K�!��5j��sD�8ƏR̗64Vkxb�M�z�,�n��k"��r'6�V[�1�v`렣�`�	v��Z��H��A/nh86C�BĈ���%��Ol��BVh���e44��	LR9��u�:�%�uc3Z��n���B,�t��̥4�ٲ� ��f�ai��giR豌8Cgd��\����m&&�l� n�Q��
K���y��]`5!
�1BҦ/Z�3��P��Ul��;����n���Mh	�-1�mi.��!2֨cm#���s�UB)(��/�ޗ>���\u�\=�:�^�΄c51��zcFNe("�$E�
J������;EN֝y��˛��Go���A����v�Dh+�_�^����T���Ar�nw�ښ!�Z�0��wh�F�b��3���V����d��݄��������vO`R��%N*���{p)��1&���e����{��-G���l�[[�~���'���{{ԃ�/�uS�d��jI�>���/a%x�w���g��qx��to����<"!�z��Z��w_l���w�D��1{�4j]O��{帑�\��Xy�XX����*�{���eq�]=����SۢWcٳ����Po�\���3[�n�7~����%�A�=�L:�<���쨛��!�T��m�@�v5�Q'$)Ѣ��^�J�!�ۊ����^��g��d���"s�C��}y��Vj�$�Ӹ�'0���[*�[�U���&ªT��VXf4n0v��麓�tl���L�ne��+��݂�'3 Tt��1����&
PW��Zpt{��F��ge��ߥ�,"w�˕�{�r�K;a���qS�؛��}�V��)�"��c�����[���+ў9�n�=��y4��{1m�uoP���J�"�Ӛ��B�Xnp��sx�1�⪽%���z0Y}�&}�
��2?)��9��ѧ^w�*`�{p�jԦn�`�1�%��,L���2����݁d0uQ�itׂ6����+���c5MY���j;�Y����.�gj1I�$ƌ��ɴ16�b�Ҧ]��ټ#]E�ZPїl�`�K�bKo���	�Zmz�ٙ	H�Љ�s����kA*��X`���F6i�����TH����c,����*�vn6�U�f]�Qƃ3���5qm����6��2�á]������y�����gP�[���╝~wn�w�u�;�肼yW�l�}1fjnճݏ�^�)��<�}�R���]g�33�u���Qڵ6�0i���5TN���Қ��cEc��䅎 ��m��C6)�����Q���
���$o�~+�2q7�TiƛޟV�h8^q_%�&<D�$I���VȂ�+g�jE����Kᴲ��r�.��W !R��C��,��]v���� �ii����tDD� yCϪ�j�Q�:�����L�t����q^T���zk˝T>�����#GB��:��B4��&T1
'�*j=��_f��8�g���� U�_¯܅�d��>�+	�>	��Gν��*o�>����n�b&
E@3bff�Y�Z<�v���9����䐚�T�uH�y���!��U���ɔl��q��B����ؠDA7��0�kn��K3�&����e�y�t��t�贌��5n۾I����\M+�h�_	�@ut�(;TSXF���,��Bwby�� �ׂ��j{��Ξ_K���*L����#�y�!:�zO����"	>�d�@�+k˔��|�$� ����ɓmxa��� QG�����J�c�x�G�|��5V��Q.ݓ��h٨z�B\ŝ��]�s���tU���5��w�X�xc뻢�6
�u�{��Q@���(8B6�FyQY;�_-u0�����F��D����7{>]�x�i���SӠ�E��%��h/��4ȿ���x�g��Lh�|'��>oh�/�"��=��R.n�nl����>��r'��·|��p(G��҅�����E��	��~�K��g��)���D�*ҩ��8h���}$���h��A�>�����0���d�eZ�}���]^v}�}�/�c�&��r[��Ml��uQ����@d,\MZ���Dnv.�G����y�J����%o�Ѱ����w�@����n�f�=`�[�+��%���������ŝ=��)6��[)\r87���/��m9&�7δ�#NȮ�;Q9���4�|>�����̘�2���|����b�5����t��ފ>.7�@�a�ZG��u�� �] Z{2���|�t��ؖ�s\n�di�g�җ^��6@��#U�y]
��]<������s�I���v����:�&�*�P���sJ�2b.X���o۾��DɃˮ�A+��w���Z�o�8�jɇ�N��q��~�۹����f�n�"��Be�G_M�`Y/EIl:}Q
HbbbJ�P��В��;��aB��ئ���̜��F.fN�Bgr�Z���z����HBf|J��>h��lNڲ��˄���tp�s������Eh�65>c�]=?�w����w=���K�keRfګe����:at��Vְ��P�kc3�`��Z�%��4G�Uw\��vS{����[^u�~�& L�]�(�<�����=���z���?����tM�q���Ua"�I�oJÙ��q��V:�޲s�� ��
]�v([9�ʰ䅢I��?����?�i`A���Ӄ~�h���H�l<|E�W��ro;3h����|Qg���>Κ�BO��!�*a$DL<L��bV���fvZ3`�;>�Xx}u�t}�6Ԑϡ�)�BK?n���ee�|E��H�`zJ������x<' �jo�(�P'ބ�v����IEM��z���@º8����#5��>�;;�׵R߸%����wG(�e=7Cڦ�3$ݸ�/�V����
�T]��n��{�Y�;`����I�:��3�B�uM�����]`̡" 3*L35��>
��핅Ӭ=��̀/{k��S���o|EQ��:ݭ���Es���^�mn�5�g0�Xs:��T�e�L�ŚG���D�t�T�:�ɓK
זgV"W�榞t�hݵ�U��<]dT��v��H���rHfm$�����[����`3�L�*L��UM�F!�ؕ��镟X���i��uB|�y�<�`������L$�if��&!LL2(y�Q��G|��QE���]�JhiO�|̞f�� b�O����=p�ogx�4�	������!�2aB������'��a��r�Z���w��x��T�ȬZ�9�K�L��V�}/p�}��[N;-`o	l'C�<�n���}~s�~c�C%���a�^m}����>�P��±{@�w&��� T1�K�5�n>&��!���P�z,I��C��#��8�V��9�%	��.�:��.	n�3�(^��f�[�f�U�U+�p�	�ܭ�ca�&0F�QJ^{f�y� ��Ɉڄ��U���V[)2P�e�Bь�[��+XF;6�G���,nLQj֥`��Tˍ.�JP��Ti��J���
��4�ƛ����)e	�"��[�(6�3P#�V�#n��nY��ZX�6&��,�K���b[*�le�a�%�I��a�A���(�J�>=�@a��N����z���8s4{�r��'y]<��?y`ˉ�����Ֆ{X��x�h7ݙ�ǜX�M\��;o����3�q�jRXL��.�5���kvn<v�ja�� �0�HiY���}w/��~:fX�L��U���i}fGcVB}}�hY��~ �d"�XGj>��cAJ���D@�2bQ�#Tс�K4C�}4��N$y�'<`��ӫ�p�`�/��+�[S&�rL$�P-,[�:�x;a,v���z~��c����ON�ߗ�B߶k�u<ɝ��7�޹�qF�-���BdQg�
�UR���15F8ݥ��3�q4��;��>$��;��ʭv�ė[���90�+#}Ҹ҅��+y{p �x2�I���f��Fw�������-t������
��:zgH��QV/x�����sa�ǈ�� ��qȥC+Z��Z����1kµ�Vy�T��
f]<(說�xm��ow�XIx�����,<d-��r@$��y����D��Ɵ2y9����,�DD��{m2(����xY��� ����*�*�#�k�Z�d
�#Ec7�� ��7��،�%"�HY�ɷ=��D����	K2Y���D���E�.Z^��We�y��=�����Og�e7�؆?q�%麂�硞�f�oU*6h>�ڄr��L�,��u(�}�
/+"��HL�O���ιB\�Թ
2UM��6v�|������#������ʚ�7*&��o��&��ƌ�\�xN�>�������Ry��O��YʾǓ�|�F�J�$�@���Mh�n^yZ8v���О<DM<,$����/c�䓳(�矵�D�}��+�����>��a"���p�}XAn��նIA],�`����n�[�`m���0
�!ǽl�9+���j}�/�}<,$XQu;��-u������	7����z��}�<�5É\�Vۛ�:'�=�ם~>�e��ߺ}.�m<'��Udj<a>�Zs$$�-��ݣ��|t3��D�/3\Y#x�3���	�}�L�'q�����	 >@3�	xl� 遻y"
"|��"�,]�1#�̐J���#V�T�@��|�=W4JY�d����x���ݡҬ����1s�Mzf��ݠ��\�c���#�r�ZG�w<n޻�,H��ǘ�3�zeY5� qV��v�C0F��qL��͛�s٦A�m�8�N���=��ϧ+D�Q��Ei��=-��,*�߫uV�s$$�v�oY�4�}�#�'�S3&�Q�'�mlN,$	�&Vw���E>�C�=.�l<'��Z���	��8����o���V�W2��6���$̶�l�ac�2�K�s��b�lG��PgGAv�8�.R|tO}�����W�H��:[��Ֆp��ث�x�G�F��?���������Y�����X*,�̟L
���8�
���a����m���պ��u̐�X*�vԿ�4�4�<CI�a����?�}�4���6�4��Z�����h��Fs��3��<�:p2�H�v�Jg�� ���]�?ƈ�xOغk��a����Ĭ(ºN��\N(r!Y�qW� �B�nI�r�'�ceE^�2����Y1Sl���x�i��ˤ@4���W�t��wih!���bbʟT���[fwq�a_zoH���g�\���TƏ�W�C�U��7�+�=�4u��/\�P��}��*����Α�o z��i���Z��?wg�7��"xN���u�v�đ;���y0�|n���}՞r}�V�>��)Ba�h�I�Be@M����@�]xX��*Sf�[e�|�:�%Ǖ�*EL̚�,��Ǿ�򢚲7v��`����<s!/k�-����PzvO�W�Rib�t�)?{/<?��Nj�䓤�%F�
��u���>2;�ٯ�ԍ�fVĬ9�MCY��P�-tX���	Od�S���Q����''6+E<̝2�L���i"�g�V����$�A��"b �33�:)��vM�Wt֊���]�F(���)�Ó	H�|->�W�+z�Bw�H��A���L�/Vj{��}a�? �*;���/kԿs�X}�����}��j9����}��//dlT(���5 ^d�o9�����8���,����򞘟JCĉ������g�@N^5���h���A��%6M-&Eme�u!H�i�)�y��iv���k!*[J)n��.��kn�]ęc�Us��b:7�I^i�⥸�;<V$	�2譴k�&Ў[c�i��޼������DtE���,
�05pK-��-�U���fwh�/2��(����!l�[e����-If+�."l�c�Ya�l%��}J��YՊ�I-X�֐�)�ݫʨm�	���r�j�V�Rq҉��4��u�;2���ӎ�ي�J�u�i^��e��ɰS�R!��oﯽo����[Rm�"d��X���+��ٴ��I�f�b��X�G+;:=;#��\O���f��k��r7b�$3.����Aq���5�d�h<!�\�~����䐒�2��S�߹V��N�8�����_�n����	8��x�|n��KD'S* ���(X7Ne=X�����Ȭnd��m,]]�z�m�_]y@��}<�[]띲d��T��b}8s�jg�%aF�{��Qb��/g���=�zO����~��s\�͗
K̂Ѱ�DnaXA���&vf�K}�B�ԟ=[�`�7�2�B�K(\�qS���ZcA�L�lh兵lŻL$��*��i130�-
,K.��{��z�ƪ.2o��Ui4T-�� V4e���ϋ*rg�B�p	�m,O�]{���x]ny(R�)	D�*$�;3ew,�?xF�V/a�˜P���3w|PW n1�+�D�u�hV7�3�����NQ��F��'���vH˃0�T8�m���w"�B�P5{h3r�=��A����[�M����^3�V4b��w�ja�w�s�XA,'9����l�s�pd9���Av�Gܬ����T�`�O����$��&)�ó��0�D��w�@�&b�Pi�ѱ�u�Y"��ɫ ��&�??u�Z��Zx��tV�;?A���eG��޳ѧ�y�����=��h��g�,�X�78�%�̅�2Vo���O�{�
#�)�+E̶���	�[�xR~:�����\vS�
��w���
0��~zi,���?��	�#ޙܗ^�Ό�M,�4�˛,Ƴ	�Lj�*����J��s��ͦ�^��R��x���������|>�ź�	�sU~fq8�9��_Kq"�z��d33%	�(ʘ�L�#M�/��|��`�a����/Kٝ��������\���x����&I�	�3���"��L�dSQK�(ם(�����
e��Q�� 9����wKtVc'�昽c���Z*`۩��i�f�N`��R�:i�{��u("��q���.r������Qu����*�x���xv�O�q;����O�h���Dڬ�Ƨ��p�"J�{"w�$V���2n}�e¾��C���R�4�������0}g.���%B�cU��s�5ϻ�����oX1��dvz�{��/�#c�':�]�O/���ެx�-Ow�l�tb���=lU���/�\V��)�}��\�E��Ш���ic��ͻ�O����٥=��}��yب�� 璔��:��K���(6�s�1b��j�����b�ѥ�wQ�cyZe<���|����k�N_W{l�QQuY�����tdM1}�&�����r��ڜN��`5�A�����螢�T�c����5T�#���}�b�X�	�!��^].����'R�>�\D��鳹ݍ|6����_{��������}0�a�&�8:�6ۼ1w�1�����Ei�R�'�J�S���S ��O	�n�%��֫�8أK���������rs�\7��Z�b���ؾ�#o�0�w����{�Iu]\$�{~x�������K/���Y���]�qVn�1�h����|>����2�F.s���r���c��ѱ�-�˻.�^�ke���Y������$���:��n�3����g�I+�B7�ˈ��[YD�ðf���v��t�D1�;����*N{��w�C�&�.!�����7.�
���+�����}T�x�����*�l����J��s��Q���,�b\X�+�#iT����u8��M7.E���<�X_t;���}�ɣ�p����9���K2����
R)SÃj�/f�E�6sM�|<T��w��!�j�����9��G^��틬{�������v�5�Y�9�x�����:�s��~ �����xl}E���)��]��9ou���B�I�1�lɦ�֍��yL��aX�s[�Ъr=6B;~�.�[��_{˦q��s�qoy��1u����!�L�ob=����$�?!��k��Sw�"\��ZsLb�MD�ĥ�����U��4�����>��2e�{�5�ۛ�Xq���f�f������;:�a`,�L���D#ț�{��wU���p�\=�޼��� �����N�'�����_W�nk�إ嘼�@�^>��ؐ�xχY�Jݡދ|y^�=/A�:Aj����]���ҭ��ew�{N���Y�^IY�y���LIE�]Kux��Ipɂo�]�ݹ�E��u����Wn���^)	�!�hiM�.���Q�L�x�4��I�઱�	<	��龧�"){�]lmڶ�L�؛�O&����[=Q{�u�m��n2��n�{�������g��<��5{���I��e�f���{&'i���N�"1V�R��,C��ڏ[��t=�T�2����6��ݜ���wN�
�Շ��b���:��1D�{��vr~�t����k�;��x�t����?=B�T����E��C�l�w�ʴ�8��QjJX[4����s���Q�K�|(�U�.+9	>�R�t ���n��˝t2[G�V��z�s��t �F�<q��nzkE���`�s!�P�kt� Ï��:O�K��D�i"�z++v+x��#�z�\I����SIb��|��(V7%�}�|�\��fa����Yl.�f�!,)��T׈c�{ej2�o��Ws} �ҥ�LJ�����讘X6l��a����u�G�n����?[��P6R���D��A
�]TULh�dl>�K���_/os���-�Y]5��������a�
��'�$��xR�^d� �|lg���Y$�u�V*�g�ûeg�B�M(Y����K++�D�L�y	�x�|�9��@@��}ʴRi���
Ƴ¸�ɬ ����J�\�ٻ��Ѕ��~B3m_�0#����h!��eGjt�ϼ��"�us6)��э�PG�@G�k*bȗp}�Y$��W���l0$�=�%��e��7�ˆ���X�:l��MC�^[v�VE!�k���#���A>&�x��V8��"֨��gP���D�X(H���VIg�I�H4��=4�)2x|(V5��M`��㙁�^W���Z��V���ћ�f�J�Ҩf�Ɩ�9f�V��flؕP�h��Xw��쌬��u3��I�3��a�c}-�
�'�z��eBl�O��q�O�=������0s��~'G�����Ù!�2Z+�]�Eh������L>�f�ӓ,vd
����`\C����9�Ӣzt_������~xȬ��C+X�,��zj0�7��H<�tEv-b霽xzty��$D�a��t�ᴡ}=\�/�����+91� f�t��]?����@lJ�I@�(J��RY�v���h�/�y5�d�ϼ?��/������;��a�p4|�돡-�ܟ�K�h �Q҈�ڃ�4�4�v7Sef�F� ��<D�LjU#�o:chq�pҝ��_z_��H|�ޤ�
RT�E�v�&F՚�:]�%ه�r�]1R; �cXWH6�5��RkUlbc�FջL��r���k�Z*Ej�v�T֩l\�MR��\:�6䲮��\mb]k-��R%��ͫ��
�McM4Հ��r�f)k�fP@l4�K4IF�9&nu��%51Xb��r֙��
�\�U���lܶ�*���R��y��f��}?��ĴS�#��^n�������cT��d�x])�R�m�: �x�\�;U��q梔ۭ۪�O,�uAH�##l`��!�G�*��A���P��SA�:m���7��!f�����a+��_�[�	Sd� �P��B��e��Ȭ:�+6d�2^t�OC�b|޷��E&+ts�L:8�M������~����C��f�S"Ѱ�}3���/�#=fC%�j�7�V'C��]�0��V��x�{��7�����I��ec����ƈ���L�:l��W�P%�S��C�Ȭk�I� "�]��\A����Y"���y�j�s0��%�^���z'�d��~�\E��\��{��s7^4�`�24I��ѽ5O��TȰZa�Ln�XA���˧f!Ǉ���4��iss��h�Qݪ�$Kef�Ƃ&���I�oS�Հ¹�l\�@��w��V/�%�� ������3	.�N�h�9����"��	]
 sXP�/���1쬨�u����S�R�&f� ��
 ݃������lڅ3��^��d�3@�-�>���q��>�<+����eX�U�/"=������wt��'�su^�1����}'k<�Z���ζ礹���x���J�9��\K�94�2>z͑���XA���y�$VH���b�\��5�u�wqK��w����\I���L劇/1�979��03�����|tTrd��Vx%K�˩�Aԏ3*��`����w~�q�O���5E�Zu�Ƴ-pX3�(��z�zN��?]6�9�vtL俎���[k7�h����db�������Ⰽ|��ߝa"�NIE�}ҦDn�mո�����8�.ڜ�@��m��EF�֒�h���M�>;��N��n�fV9j�!D���I���	,��)��xr�9%���-����W/��-y�y��^-�s<9��6���}'/����h��E�|�b��d��u�܄��9	:������Fa�����i4T}|=�+&��O3+&�Ry ��fN;C����}����]tf����� S��{��ԗ�#�2HZ��vR	(�VUe�K���v���� �Ꙩ�n]�IN��r>���<��C�[�PZ���ꚩ�?�ח�̚���*�\  �Y�r�3dGO3L��0��eI��11L˫(W�;p�����P4����<)��E4rHK�	Y&�<h�ӛ�%���]Z
��:����=���Ѱ��0�!	g{��<h���KY&�x���X*�$��GLL(t�F�0�Y��Bm����H��9.�.�t+��q�K'��s֥�v��GW,��(W�_M4�)>�����yEs78�;=?��Y��N���yn�3jŇ�y��XQb�qQ����e�e[�0u�����쬘YBy����S�^P����ރu����inv�-���V
<^z�Ec~L~_�dwYZx�P����d��q���bfQ
S��L�`�\�����c���J\��4�)�ǋ$Vw��|$���-X*�ࡠ��C�4����݁#B��$ꬵn�I��z��y[����W��,�(�Oh�}vQh����ꘛ�X������q�66܄��QW5��-� �Xc����&��]ix�6Eè�C�O�U>#�	�}�h���qέ#YBX��[?�vO�
��7B��c��Jw{��]H�F�ˋH0�03w�xw6$��"ࡱ�
L�ۮvRm�fP���l��&��ω @�����n��8�a�O4�*��$V6L^*�Ag��T�ɱ�Hq��O�\����v��} r�9�P������/^I�$�	Ƴ���_sɧ��>�M6�*.4|9����({�=�AD)u"�jj�p���T�K��&s
�f��&v���-(y;�����y92)p.��U"��L���_Os�9����x�cC��s782;��p�P��wt��H�C���KՐX�s3Ь�Y<�:�C^�wEp�o;��o�nWک��I\��_;�U�D>�Ow7S�=���������c���T2�]���L	ȇ�O�D=�^N~�]=os�ӯ%)�.�\-�I��-�B�q,�YsU�<K���\հ�b:�a����*�.e�m���"!u��SL�T�N�e�T�8R�$��@�^j;:�� *R��5�,rc8��m-�Qѣ)�q6l̴�5�ڣ�k(@X*�Yek͘aJ.�V��m�2�����f.��Z�.�U� CF���L6ю7���^�J�[�8������؄�w�.�v��z?���D��7���e)״�S��bk$K��hDΤ�F͚�+F�/�&���gS^[�`�����ͭ{-�8�+r������i�����vb���w��]��gmc
h�Z�m�k�����5`F�O.LKΒ/��RY��*dV5���=~LW'��*���(Zx�W����@�U�xLq<�O>䎗!�|'�o�h�r�0�X�1x��>��R�O�����Tnu��<H�҄���VAb�fz�a'$���ǣ{��P7�ێ�XIg�����iWC�5N�������I;'_}���Y����xʘ�ucYɗ;2�ww��*Ů�%�^S̨x�k$VP�VaV(NIΐ e���- ҄��4*�ǌ V7%�N�``��3m�j:6��v-h!��]aٛYY�R�3�dGRV�n�ϡ��']��5SC�̪�I��Et����>ecՐX�Y��\�70	��[�z�xo
�(|�D�R�LL����fW�K�[_d��vE�tGm:�@{��ϸ� $1m��2�zG�h������La��zτ��%��8�MWZ���bR���&��=�$�������}k5��]r/'����N�L�5q��nظ�mTE!�&N��@�К�o�eF�̧��x���ug$�:!ib�#U0◉D���1\A��WSҰ�Y�afaX(�H�h�ef��ȸ��	�;_�4/���p:���w�O>��b%9�zk�&�S����9�Y���@K�t����u�؝;�����"H�z�@����l�ҏ��9$2Q��b�ER�;��,��+�s���-���U��"q^s������5���g��4�-3���̳b>��z7D�]�U1 �m<(��+	,_S,(Vxu��=s%��2/�g�d\A��ϟ�-%���q?��_������$��O�ʸPi�Օ.,���g$��&���}�w�<ĸ����<̮ ZI�]sՋ�x��L�	;�EQ�|6jy	�D؂�E���@#8.j�B䡼�32=/�	ү�}�Ͻ�x!�9��D`��!.� %Ɉi���	D�j��v��_�ɪ2�P�!�L�S�y�i56gԴ�9��E"��0-^�lDmiP}�s%�!�A�/l]��Y����=F�!C��:D�������y|��������֮��ty̓��X��tJ��xY����KT�+(VjH\��u�.���
�W`n��^4H�q<1����;�q?��N�p��~� Z4to*�Ag���d}�H��`HbRB`!3�� �$lg���-�KmR��Բ���E��Ąh5%-���-�+��S�svn�ս|c�tO��v�+$�������b̐�X�$�4𗿾��s�?O��Y��q���a"����zÙ.v,��OD�O��<X�,��Xs!� e��}=����A�����o_O���fY�Oמzi97:@�����x��=w"~?�<��l���p��a<�t^W��i�E�vO�a"�O�[�Y��$�HGšx�W�h'�pfx#|PF��b��E��DCĿl�r����$!�/N�'�p��v���s���Ns��`-�;�*6E��:�o��UC���5������ї}�~��0�Qv&'K�J�����w�~ع������xOl���
Dw*�\��"��'��B�g�������G!`�xY�Y�/�B��\�"i�&n��m��*�i �#j���,�W-�$��T;��{ޅ��������hZx};�5�����1:�K<)���\����x�X��<i"Ѿ��D��P����U��'���u��ܗ�p�$��O��z��}+	�}SxU��rp�9���g��SG�5�39l����+�i��P����A�!rC!6{g��^4�ڞ�g��fC�ǔDü'�(rfb���M��	X����ZP���w�kIv�酅s1��@�
������G'��S��N<�đ�K�kg��Ta���6�� :��Bᴑ<osՐX�I�P��Y��*Ȗ�������f�I���w.�5��1��]�v��>�t�甫R�}��ώm�
2l�������P�&�`��������>[;}3��ds�v�$�o�w�o��Yl��QY��"�x������t��:hg:�I���2�n���}�w`i������f?�}�ﬖŏrukun��v``�s.�N�W�nЃ�y���"te�������]�N����O�C��wޖ�f�=���� ��]��vPNۺ6�W9�ٮ�����}_��ʂV�tI��p�z��蚦�jH*kdL�s�KN��Q��k[�գb��\[���5=��Vs�5���/r+f��������(|e,�ۛ7�^�Ҋ�>��Xu��_ck�2�̍��U�w!Mݞ�oY��d�P�j��ܜ�/Nv�B�Yد�M=ז�)!4���|�9�K��"`�����BY޲O(Ϥ��b�u��9���o`;f�v'����ن7�͍�i���x��f�E�О����mq��)��['NI&�o��[�r:�Zq{,��i�gC1�4�zٹ�p�z�ɹ�֜�\˵Uq���ޛ�W��I�y:PP��<��v�I��bw&N5hŉUr�=\��;���nx��I��o��Y�>�4�3���a�F%\6_ixDv�CG�I&�.��sj��s��I�|{wi�r�ɔF��ܘ�J��ѢxN����}���ݒ�]�T�Tۃ�VIw..o\b��/{��]T޵�b`,�$��8{a�n��@��e�Ӣ^��qt��{��({w���}�__��O ֝N��s�o)t*��3��{���,c��#xr��$؉"�(J	G��b+����J&���,�Ӭ4�(�rj�#�9΃�rl�)u���[-�A[�����
�o)bD�m�r�᥈�l6`C\��4�`���ܲ�it�]��ޭ X�f��jYqv-���!�5�)6`@�Z��Ѥ���U�q�E֎�yAĲ��).��n�a[+��ґL�-��q�fq4M��1m�-m��Zn��mM4�1щ�š(A��j����n#�;F$�[�R,3�\����Ӄ���6�l
��lh���`u�Y�M,":��]�	ee�릪��k,XB���Mm�+LXp�u%��t%1su���- J4�Ίb�F$�A)���AYH�m!��b�a[��mb�5��֤GEfr�Z�K��u����LP��5���n�Ld���f�`Y��i�CJ��@^�+�U..l*L�)��P))4nѢ&�%f��\�rU��Ha)��n�l�]X��C1�3&��)��Ż�sf+[����^8�LF�
����ãqN]w4�u`�3-6���BY�g����N.e5�Aإ��[���t^-	��0��+�K�Ժ�Æ^&�,�Z���A՚#R��oYN񌮬CA�sTv�ї%!)Y�����35:�
cq]J
�-�wRm+�\�+��e�1\\-!t9�ؑP��k�+KR�r�a��1�l���؃H�Q!x5��]�ne�ے��l�A��A!��F�V�*Q�����)�hEZ�5���5m.��3^k�݅ 퀕�$v�l���e�E +	n��#x�jl%4#�c���-ڴ��(D�M�`�*�ln�-��h�@�
=���-:��-J��YfB�ji�-��Ŕ�vnֱj��1�$׋2�gGX'Tw\�P�tpF5+t�5\��`��.�R�m/5ڒ�F�M\%+�!��#K�tv��bX�Ce�l����z�;L�R�^]@��:�b�jFmVi�`�m��[�1Q�T�&�����
J��$)i�6c������ބ���׼��[Sz��6��~ �E��V�.G��y��)'帷�ow��g����sY�G�ՂQ�t���y� O7A���\ۋ����Ǳu~\��T���.�fl�Њ�|���˷�.4�g��^�[Σc]}4�xDz}��%����࣊z�i�2�Xf�^>�cM36��<���^��YJ��G�_z���f�܂����Ŵ��"1V<��@;�q�6�f�+u0���&K�g�۟��)6�ϵ�&�nK�]c�v��ΥrРC�7A��pk]�*�Z��{/L�-Ќ�[�j��75箑݃x��-�`�ލ�������<�Zwѽ�3��~�Z�'Ϩ�q��Y��j�yt��VL��5*fٶ0�^��Q�ʱ�]�Q�f1Y����tf�$�R(�a��F�Ⱥ<��o��{n�ub	o"6F�Ëz1o�ɧ_�	�ǩ�5��=��sY3��$�1�tw]����Yb:�+��l�&]x�9�(�<�܀�N����)��n��Xq
{8D!��G�z�{���]F_w��)VE�~��j�ۇ-���kV
A!J�tx"�[��7��Û)0[�)Ù���`�q~3t�d��v�O��?H/���A��^�M>��w;]�;��=�r���מp�O��s-��^Iw�Y.[99����N���fR�V�(��ôJ٩�1����1�+���T���6T�%��AH&��Z`���*��p�ܸ�����i�9�mM
�դ3ͧ,��v��R-ne\�f	V�b�VB�8j���ɦ�&]l�:��X".��h6��ƕJ�\D$�-�݈q)p�x�!�1�5v��l2�lv�` �$m����,�MR�#U���4�M��8�3+jl�c��j�=��Ő�qن������f�e�B�t!7�)�5�P���<�����/oQ�H��xt�{�y+�K9���3�������-,!���JJ�u��1r;8��,uj)X[���K�R�
�<��HHFw�F�79�c����ts��:�.���	�=�L�O����r�d��):���x���x��"!�fEcY�d�b�����$�E#��δ�iC��ɬ$|������i@��1��O~���ћ1ٽs��H��"p�X�1y5b�f�`Ii�G� �m$]�U�X�Y	ʅ	��A.��bbaY�L���gd,>��z�P�6�:]YE��fM3�s29!�>'v:��-��C:y�R�1���g��v]h�x�a[��+�4^�T����|7�5����J�G})�rH�%���e�B�`�%i�n�V�v�Gh���X.톚�U���� =�a٬h\�i�f]q&��w�M%�O��xc[���$.BZ�ƖtTr��#��%Vg_�����:���ݓk���+�^nw{`Q��J�h�Ieʰ�=�'ѫ��W�-����DQ�����G�Ŏ�a�77wTx��y�旴�U"0��FN)��o��,�0o�^����y[��|e�֣qs1��1ν�!�*�ٙ��I�!�+쫊�P�>��N���	�=�M��r  ����k~�Mغ�\��F��(��<Ldb��.N FŊ:w�q���#²d�A��u32ҡJ:X���b}�-�9��~�> ҅�g|��X�s3�g3.�o���|Lzt&�ϭkY�[�9��5�(��*�,_rI��	�/�B��̾��i}g%6�GM�����p��Pn���* ��Z�XCEf3XXM+��cF�ێ�.a��W���w�4�+V7�g4^�tN-�i�͊�I��T���2�ibު� �xSj_����0K�/3
��\g�&��f8f����lt��M</���SQb�"�g&c���u�j��O!ɒS��/2�1Z(4�:cڝ`�H�gt� 슩� H�VDLǗZ��tZ��%-0iA����U��o�&��Qbh(�gкJ�q0;�nM�LrV��,�����w����\Dʁya��tn��^��������Λ-#�a�������RJ����oa�8�%�r�B�ƚ��j⦳>�|O��u�HdJ'��*�Cx�#��D�
�D��
/�r� �����zh4R-�؜ V6NN=`���.v��o���:�m<'�Z��w�-2 ��+,_VT,(V{�.�!��-���F��K�$���ة��I�P�a�� �Sg�B]5��Y�]-+�V+7T��f�c0.?�zy�����l��%�OL�[��* ����z]t;tW~��I����N�k$Q��W���o��t�-ZxX+�}%(@���S"��>�����θ`A�����<�
���Ǭ3�5X�k�ʔ8D�D�L�̧X6E޽a%���#��e���Oo�\(�������/ʓ� E�P3����9�9HD�����x�|6��MX���C�'X5��.�CF'��M�I)T�~�Cƻ���O��E��X�[�l)�&Xl��tʾ��ݷ��f�g��0����9���� a�c黗�t|��9vڜ33F)�r�E�w&���As�$���`3FU�=F�7z^�b5?����o��/�i��h� A.���@90��u����U���re��]�O!q&�'��E��/�>���'�B�.&C�٥�Q�(6�ެ��A�����5f�f���cϧ� �;{�vb��ж�e�|Lzv{Ӿl�s��6��$�|d>y�$7/������c�q5���^�7�b�V!mU'�?��=�K�'�d�%&���GC���c�k�X�a���``�i�gu�f�Urݝru���#��3���?Nb�rd�!� CX���Wi�_�w���D��,�J�0�\�Wx@��� ����k��4��~�����XAg3s��Ba=�b�	��_�ȗ�f�v*�xLq7�� �����B Z8WOc�A�������X��5���%�/(���-Ѩ�i�5������#gL�]L&qO��'��iV6��}V��FY9o;g3�a$9<
DZ�D\��MaK�
̒�`z�b6V�e�قW,��f3�pQq9��M��ͮζ;Tx�5�6��͘�LG�p����:��%a���ml�际a5�Z��r�6a���݋��k��fԁ0�э5�3X��+��"+V�PY�c�ƥ5��n�*��3���`0ġ5tV��3M�"4����(�v��6�`����6HǾԤ�y�G�.K>[����.�w׷�.��-����nR6ܜZ�7w|P\��.�fN'�{�O�l%��u(bn]�%������j����p`c�\^�ke��[��7W�{��8pc�h��n��e��Bϰ��.��<YD��(�6O�X�̗:@�B�|5�'x��xa���* $SC�1�������5�&B�!�u�w���&�&�:����U�$��  -�X'����ث��l���O�}ߏ^��#��
-��K�&�^��,抇�ǣX�Q���� $�D�+��>�H�{�r��E<����c��K��@�X�O��h�n�bO�k�lBlcC(���d��ߒ��`���-�ޘ�E�t�S�
u2�;��!�3d| ����DBBbaJ.u[�dl]K�acY������35����MH=�o�~�p���ۙR�f������+({3�5���_3~�9%�a���ib�����h�}ü��ǅNQ.����0�`��5g�`P_���u�9�9�	>$�DlQ�>6�������6��#޲<H�"`��I�[!�kFj��^��5���k�}�;˺N��s�g��6��(U���8w�1�dP=�8p�i�[��40��O<��~����ש���k(]��	!�Y��ً�V6(��+q��X�gea̅�'���/A�e��Y��o^���|M�
,��X��䛓�]8�u���@�h�U��τ�Q�/*!<D��3#��2u� +{��q�E��a"����ɬ�7'��/>w��\Q�:}�LByA2�&%餱x�%�$[����:`CFǷ��Ri�c���E9�Y�I���tm����e�@��mbbW/؅`9Jds3.���	q\\��� �+/F�̐F�t�����ߎ���Yu�+
,�2���n�;x�x��w�'����M4c�:���c��1��g2�(@�Ş����SsҰ�Y�>J߶k�u� �	'W���V�6�T��g�G�d���W��,��������>$a�oE�N/k��L�e��}��Ƙ`Z+��U�����w�Z��}�1�2T `Ks�lm���B,�8��3N��n���O]f�e�s�_�	��{�{�玟�\��z}��=�m��xO�4�y�|�h>�'+�����mz��I��鋄��!b +�ĉBy(�>�9�[��	���i���[�X�j>.��aE��&\ d+u�r�'���������E�UߌO�7�8���ώL��p�G���:��xQ�VX��T�(Vx��gP|�h�X�sC�H�J�U�]T��u�Cq�&�U,W�k,�J,��?��C��w��[����\(O�Q�	,�<�c�9b���?3s�0.>�F�=h����X�R�\��"]D�̺���I��+9��X�!x�H��Ҵqi����T5
�2%a��\�ib�����*%�bf&	��i4T\?dŐ+3'�Q��8 �X���c�֍����XId�/�to!t)�f�n��O�I/�X=��g�\(O���XQg�7�覂�J���FT�ܤ8��0��{Z�ىm)8BK�L�S�1�<�C�d1��������A�Z|�Fm�S��Ϫ��\Ъ_��d�U����2����KӜ��k���l��}	���8yi"�ť+UR^�ծ�ۑ7��]�0_{��cF1r>�ʇ!�`4���`���EFˬ�93s;*@��⸃E��OB��f��ٿ=`�s��O�'W�o�a��m
WX����m�ͷV�� m� ���\�6]�2�� !.�[�P򜉁<��������x[����K
�2&����Q\��B0#�Y�O�0�m<'Wk��!�Z^ɉ*�,^��90˒P��u�}���,$���U�M̹:�t0�4V{�;�fH��X�U��ӆ����Ă���rc�,N���=�ZA��?���g=;<��� 4ZE�JfX�.d%�C����+I>��[�~�i0T,�ț Vs0˙  ,�w�q;=?���^�cu�2��?k�z�Kܙ? 2��+��:��TȎ^���Id�DX���Xp�^��`���8�LO��{��c��H���ˆ𗄤Jf�i|�5����G+�ݖ����Y$(�d	��óe�f�.�7W�����WB씮����v��z�pWB��
k���Ť�Q�P��ą��Zɵ��l�EΚ`6+���,�.�4E��۔Z��S`rQ�f�)�h/V˹�(܄4N�]q�K�WCR"��vDm�,ֆ��T���<]�j�"-�Ҝ.�hT�͍��.��5k��mA��rld�h6��X�9=�}����:�%�|`5���'����Ve�����{F���(���d̰,�o9�=�P>�V�E�+�+�]�S��-� 苈Qq���q��3K�6�@b�}l8g���<�y�c�j��'��gbl�X�}xU�K<d>x~I!$.O
:{����bt'���	�DDʱ�e�^g&C.a|�;8��GC�(�¾Ͻ4�X��3&l���h��_9
nhD��""J�x���c�Սg�M�XQ��А��X?����iC�]�`�i.o	a�����̡Y%�$� �Ft*��i4R-�Ȝ V1^b��d�8� Kqc�:]|6�(�}�B��y�Hyx��z�KT�+VW3t!	�����h�7�3x���xY~�T�X������{,ҍ�p�� ]M\��2Y�c*ܡ���m����YX�A�Q��^��Yo[О��^�4l�-��bzs��:𝟏�Lf)V5�}7�s$q�v<,w��1=:?o��sk�sb.����c��; ��� KYs$A�Q(f��|;Y A�>�R�۵1�ȍ��,�.EOL�GTyQHܮ��>���֜�Pǽ+���yo�C�Jc�]W㛬{ޣa:�l~ I�����{�����L.�3W��4 �*0�_ӖSI����LP�b30�2]p�C!x��")���f �R��˫IFg����Fdǅd�����xϧx���_(XAg�珁/�c��Wk������>� �t%���:@�h�z�Ag���'V5��rt +u���Zx�|.��@��]u��'�O�e�u�_��'�}M����i�do|��X���&(Vs�s��/�� ���..�gXB���YYv��+qMnȋu��a����@�/o{��b�7f�o=;=���<9�I�|°����%rHMɏ���Za��^µe<;�qCByR�1$,$����b��73��E�;�t�h��8���ω��B��!p B������f݁��W'_����D�$�v �ZD`'"����2�A)��Y���-St+�O3�l^����|�O����l���|�=rd��C��-�=6���T�r�L�Դ�v�aֻO��Ͱy���O����B�Rn���1��p��ۑ.9�7����11$�e�Y��3c^��W:a�\up݋v'�ˉ��]���У$����^�j;�(���׾�J��Hm�'T��'����%se��d��c�m�˱v4�I��	����v�K?�}��@��Z�W�{b�ow8A{�F 4��E�s�VKw(�z�LSS/�;B-�c��f�n�0rnOt��vts�R�˖.Q=JP췪&6-�&{�SD�ֺ�ż�-O����6/K�f�8�6�L��nGVũx��2�z���z�F%��]+�}��3���}�U�i2V����yx�8���D;���������U�Zq��7_L�g/�Zd�qk���ﾏ������9-cW���i�9dN�'��������&�,o{\�jk#�N��L,Jv����1{1�n����x�s H0p�Q��+�%o��?s7�5>v��xW;M	�}�����ݝ͏]�L�e%���hlL/�䲥�WSwW�\e�C��/(��3�ȳG�Xp崔_�8���b�ҹ�p���/�+�p[�tڡ�uX�O��J�@Wy����r幤��ˇLX����#.�I(w՜'�gY�X��ͱ{������]��3q�&'���X�V�ϸ����uO����S��t��9�7�Ow���JY����6���.=��bξz�̀&#C���6�#F=�w;����7q��a�'qp��a�k2?`�vsK�Y�x!&E�}|N='�U[��Ve���^^}��q0��!��s�.���1җ�Od���/�n�^ѐ�~�R�D��Vm{F�x�U�:���x��H��fl��s���3+$��eK�lm��Tl�!�*h��ؤ�����.�p��}ʨ���Ор]*��1�}�H�k~�􂆌b��V���w*����l�Mg��=|D끌�r���sgx�y�,�w���]�T��s��۪MFu�D����Z���y�
�4-��[����� ؗyR��q���X�@p�a[��]���B�zJ0�\`���f/n4��sz`ɔ�7���o��������n���<ׯ��d�v�ݭ�{�'h�n�������o��O�~[���
Uǳ��#ω���·����e���{<w��P{�<F,�䯯��a�m�3^s���S����i����s�� �ww��˗g>^r̅���gd7�G��5y:wzu�}�w���p����-k�9��pu�E���|�.��o}��-0͍�tdw�@�a��C���4OL��: 7r´l�]�磚�����{��{w5���ݹ��j~�tF��?���9�h��C~+CBy��j�y�6셚ɇ�oT�p`P�.�*S[TTx�/��QhnЗ��(Cti;N�:�k�:IFQF�ܙ�"6�j���2�Y;g'j��H>:Q	9M�#��4D����q�B ~�D��B!D�ɤ?2�HH@�[���x��K��E�9�Y�̹�0�>;��[H�>�;�K�̩Q*^fJ�xofa,�̑�����M�M�����QX/|s5n��Ա��
�@:M��\��mʰ��%�hi�Z2�м\j��Be�G]O�[l�e*x�^�$J�	���.��~����E	�ef���	h�o/�:⏆���7Ȕ�d �2Rf~c�1��p�%(c�Z1;����OS.�k<,��zÙ��@�/���}t ��'y��Z@���Ob����0, ���.���h�O��l�X�8�D9IL�y��+����������Z6���Ma����[���\`�x��W��������(f�����>�y��	��I2��1�1k�
�IU�՘�WӦ{��i0��o�v/L�T�i��+��t04h���Oo�c8'�&+n��n���{�Q��h�����4�	i��g������i���\�@��B�K(Wy����s%� 0���<iBш���x�zɅ�Y�>���ޡ�M44������H::`q��tq��fu�u`<%śZ�ر�����X:��;�+�v.�o	�:~���%�>��U���#�w�L[� q���N��I���˭��V�N;1�aX�Ne�$��HHl�i�|�SF���VAb�y����`�@s�=?�<���*���m���c�u�b�YB��𦃙.gBB5Ջzz'��F�=X����p|�u�!��b]�|�� �H�G���s֐h�y얱�e�V
�ܠ�!�"���}��ǧd��>�6B�h8.̪g,TY�8@�\̆�����{�p�i��2+�
�s&�����
W��fJ�=��,T=WȾ͜o#����y�$�,H�f��SO�>�"݃���bd&�O��>�����x�D�8�/ɕ��L�l�\�� �+`j��X��E5���qJ6ZR�L�DCĖ�tlK"�,��n���\�jcA��4��6z� �c��Vab�퐠��̡m�LF%��]j갎]t�"Whe�ĵ������M�k{ �B�t�֘���X�6a�0ҦV�[1��SSG"7 `u�qhLۚ�fHK+v �85�%��4̔�����x�ܚ/��v�]Lg%�6u㼋tHq�-�A��*�a"��PQ����t��y���;y�|&�W��~1�@���f�)i)�4�WM��.��J��c[iY�#�,����7:���a�[���e����ׄ�Q�Q�VIe
~���3s���Ef�WztON?���v�l���z�D�x�zɅ�̹(���O���*g�V+(��Yb�ܝ	�cY�߷��T3\�|cӲ??��r�/Fd͐r@��a36{���x��i��g�p�YN�fD�L��Y�����zW-<?U�����˨�+$��!��^��i='g���9�
5�n�s���p�~�V(,��#�c�@
�/��҅��a����B�d�ۚ=��x"�3w(@�Z��3b°l��;f�Zhv2j�b��D��ߧ���/V��Uׅ\\�p�jwq*�,�&�S9b�3"y���  e�Bѣ���|Z'��u55X��	���x���y���#d�G�y�J,6�Xo	�J��UM2��uv��amQ^}�J�"C7�����>��.	���W�fz�b�A4��F����b������p���7Yz�	=^��[���ov�%`�3����$��Cx�`�oea�{�X(���B��0����O��4�<Ƞ�hO$<�/M&�×��d
ƌ���S̛��Za��./��E��VIb���;�]���].U�	?}$������}�r����.+ ���L�˜fF,oy�H���zw'ĉ@�L̕��g��F!X�x��ڄ���� �xSҬ�Y���'^����u����`ܱ�V!�y[KK*8�vVgK�L��I�f��(���p �����0fqk-�I螝�߻�q,^�c͐+3
���@� ^~'g��������D�����ݔY���+,^g�U�̹'!�Z|g]r����2\VAe
ro7�O�9��O����z�kl�(pfb4�h�Oe��g��F!Xܛ�vΏߎ·j{ڞhct���o�����6
�T$K�Q�Δ���4�z��0�vC;��-��gӕq��/�W�f���kш�#���JwD�FxC�w��E�=r��#4��ɴtm��B9n-ʙ���CQ��"@��B�ݵVI��S��qY�,�^��]�]1[��=xD�NO�� ��w��u�xO��E4)�c�+9���HS��p���?|n�-u[P�ZO~m����Ė/�2���d�� �\@����X/�32\XAg�̔R�ck��x���.��U�/M�����.!ˮ�V����k<��}n:B^�Ϟ�������g8T'�ߞl�Xљ8���ω��G��!	!Ѵ�t�� �xi�O��Q�ֲܳ�I��οy:��I�q�E㻮`\I�
�+馒�"{�y���zvv4I�
@���O�Rm�<%�?�A��yi9��1.�Ĝ�}��� B�P.�\H����r���>�px� ��bd���_2O�]�����|���x}~ȋ V{%�4ȳ��>ш
��H`�Jey��	`��٘� ��cPC�{�F��3C�P�<(����s@֎ɯ{1y4:��5�V�s3WܨEաT(I݆���j���f�Xm���D�%��DO����
\4�x�������X��\3���#r�ҿ��8�I'��ooО��vO�y�=�P�3%��%a����qY|�۰L�!�*]}�P4���XIe
�s馂�'$ůgS{Slh<��:^0��!��������q�SQ�c2P������z��/s���z��f�1<@�b?~�V
<=�d:���D]��������EB�J�E�~�y��mWe�"���~'g;7�x�g&nJ��L�=j���/����������C!0`B9�	܈����iB�UZ�G¡]�/�56�|�p믾+EI�߾�xt~;'�O�M�U�.��G7�Ig&\�@��tN�-���`���A��g&\������+�4_	��*�>K�C�3+	�}Y�*��rc����i&�T�*g,TY��4���>Wd{�.B�x*A�b��:Y^Gu
ΙDI��0����-��G��GWt�鮟 Eο���^��w����\X���3iA`��hQq�&6)rr�4�TmC�8����f2ۜT�[He�ԛ7���쒼�b1���h9Xr-�m]wBkt{	�c�h.%�.%nd�l�7��%A��0�%F��R�]�-I��`�9�LF؀\��&�v�m�UHnEn���rMZ��F��j5��J*�����0���1����0a��g�Η�*�}�^O�_^y\����b?*��x1D�^�;읞�t�3�r=� ��[&{t赩��y�ɝ���o�8I�#xR�	rƲZ��:͘G]����sQ�l���ˊ�};r�{�wb�M�4.g����5
Ƴ�ɜ°���"�̹�Ba ��Zxu��V��{�J��w"�����aE��VE.K���&�ű��F����RY�����Vt��R�5���O�}�{>����1���\A��=R��YG�7�X��˓@�ewG;� ���L������ŞBۓ@W?�O�s�s8K}��|LwH+�&s
�9 nt!�b�{�h������;�y��)���P5[�D,(��2�N��q'�g���x[�6@�h��z�Ig�3�}��D;CL�O0D�%�$W:)\ll�p6�1m@�T�u�⭎��	��@෮��k���Uu����GN� �|,�T�$VQ?Nb�e΀`BE��FoK��4���]21��`e�r���?o<��鉭�[���*��d#3#H�`�����*�w%�`��� {��c"y{5,��vCi?��ϥ^E���w\��L�. ��۾^nW8ǽ�y(���˶fn�\Of�jL���M����$z�g�{�Ȳ�1�H��6D9l����B�V:���D��&Q1;ʑ�dZ8���VaV(O��!aG2\� @6��ٽ禓E�lvDى�������`VҬ��c���@HaY;�r�\6�.��U��*3=R�H��\�`�@0���w*�P�>�:I�D,��U����>~�c�=̗$�@	����F���X/|Gy�g㟎����{���Ж�ˍ�l#���t­�$c�L�-.�.q�B���E�����	�:�S���a.f�AY��g�����X�ì��V(O��"9��@ B\|ib����I��m�<�M�WF
����<:��}%! Q���G(u�iB��ɬ �P�=R��p��<���O��>]i���"ۨ9բ��_dz]a%�)���?*W�O�v���}9�de8��ڼ �MM�$�<�Ǆ.�����g�@� �b����4���.��WfN�DÃ��hƗ/�ì("�ם��m�xaA�q���ԓ�����7T�gL��{�C��ov�v���7�X'ĀAdQ
�T�4������v~?���^鬩��e�X��2�P$@�1b��q\A����Xⲋ�Y�V(�s;�;z-�q&�/��Y�%����"e騱xW�6@�\�s��!�+���A�����A�i�5˹�d�~ �%
!���&s)3.�Xؙ�l���,t6�m��TLGPlC�p*tt/Q�V��f�-$ʞ�X/��#��	,�e^x�L�;	! �Q��O��:@�bΨu
|	�y&fJ�x��
�P��Ns�a��Y�U���T�
��L,�*��c�C B�k)���n-A���|'�D�}������̉�]"Keӌ���Q\)4�譾�~9��G�'c�.�������,�L.	�c��-��J>��U�e�0�~͟qG�I���f'��G�ە18vW�ӝ� �p<НL  �]�/0�����L�H��8�a]`��1}�Ȃn�;O+#p�jeP���o3� &;��ѵ�tfj��N��&�Oњ�hy)ec}�h�� uT�|H��vŭ���a�^�!�̏31o~�s(��s%��.{���S��ᵷ�Z�������% �#\e�&s�5ٱ�F�6*⫶�)"ltx��gl�a�~�9�w�]�ط8Vi�M�}ݿ{��s�����l7x��^�f;��>]g~f �J��T�3*dF��p��J�C`��/�s����bʿ}�X����?{��|o?:���j�uY�}�_eE�����u̗3Z�p 7~z�>��:>e���NL���2�J""$�߀
,��һ��^篧ϓs^S��2�C�!�ǽ}���ٽ?}	V
�1�vɕu�Y8�<˔�w{�:6m��7?Kt]m��v^��_v*�dm����YѦ4��=L[�aI�}L�r�񛌅bieL�j�;�w�X�7�J�b��r{t��S��P4��ht�Jg��b1zo��h��'s�=�	�9���G�^���۱�Q�SףwD��*�I-���9��S��	�Q2��O3��޽u�h�N��76On���2�Gq�.����|}7^�܏1�$�O��J���?V��_��Z{�8݃��Gf�<;���&>��]�x��Y��[W�.�ȗ��"�Ų" %��@ڀ������tC�ק!� ��p��1�f;��)�~����Y��p�RNQ�]5-qbj��\䡻��������w`�n�AiJ��]�C{���*7�Y��V�<t쳢�����q[�x���(Qo�e�8���~��ud�Y�S���������]�τ�\�Y��©��V��y�5,�7�3ǒy0�/6�ek�Y��<��2]z�Z켥[s]sq�K�����E�cT��0���q\��9ݾ=��y���.Wj�WU=.軈��T�?r�ӗ�n*d���H���w�y��R2+�Ž�jN3����'6#l�r�"�`�2+��1���=ǭRs�lY�'��ͧj.)�s�l�������c�S]fC�4Ą�����v����ML�]+��մ�:֭�$�j$-��x/h���}�0%�'��i\�j �1����o�]tUɾ.�e
jM亵��ؚ��굋Zf�����΃l�cg{��0}رm��ڸ�׎8�h�������5qNo8�Q�8��xЈKzn����<��}��X��[(�Vmf�f[,��4��U�+n��BjK�k`K�Ɛ��Vc-[1�XB�a4p�N8gS]��$�X��f��I�K2j�W2(]���a\�\���mJ�st����[��֖�9&���k��hC7gT�U�2Ų�0+A��96S[)�*ˮ�5�7!��Ni�!����Ktv�xnIVdr��p�L�&���Ω*1�p���3B�¸b��<�v��V�$K��`1�\[*&�j�eteuL��eD�8�t�h��l1,��Y5��)-8(�5]���f0]2+1q����E��+�J�kFgK�B4�ռ9�����6.&+�5i�����z�(;�d�e�� :V+c�v���$�J�S�JT�ҳ
6Kǋ���tr`�����;��wfؐ�3�� �f��RmV��c�ؗcS(�fՇ �K.�) K�CcJ9t8�d`����f�Ze���%�ڈ5! F�SJ�LZ�`��F���+6lʗR-��8��U���1^����p�!I��kE٨\��v�.��mB[�Mr\��4ز��.��f�
4��YR��5��K��ж���r�!�fJ^Xj�����Z�,�D�B�T�HGx8!-%Ń"ݥ��m4�3��L�T�<�M��)-^1��Y�Vjһ�A$�[t��L��M�y�!f�v�� �A5n&V��5�ֹÔ�Eu��%��)Jˮ�u���^��l�˯37L�lq!��L�6�C�3�LF]pb������h��s�al���,���&#��u��n@;f��MF��qv�%:����Y�Q��&�n8.�33�]�\����)�G\V5�h� 6��,e�-���$شaxZ�r4��n32�-�\� &B)�qW��3mm��q.YmLY`�1��PsmM�YMs��"Rj��
F�mc�BV�LB�X�e+�0�7-��b���Sr�,[j;FU&(f6�#�5���2]1ֲ6�h�.�bŌ	����%��y�5��zv�$��Q�dD�^�*o��S�h���� ����̻�a>ڼ�1�,~9�g��tD������/{�l'��Zv	�&�`~�D�n�=�Ş�Ǖ�-�����/�j��D�M����@�M{2���{؊�';���b~���$�n]�֭�p�j%?}Y������pE�'4�yi{��\�:6H��_�z=���w�NB(�T��QUf����p��y�����M-�������*/m�;�p��K�
󲌻�x��gh�k÷���=�C���dM��ްKC���4G;{ֺ{�n��N��K�������{z�G��� ��v�v�U\�GMXq���z���!��<����*�y�brR���{�ۻ��]{}��r�sW�:���[��
<Z�'ݐg�D�;�ۇN�AfOg��ʖ�[8�Ev�4r��-ߛ&?W��U�ߪ4��k��#
n��W�� �L6�dR�_QG�8t�O@��[;�>v����m��i�$������.ź�L�}�����~���K�0I�&d��$<aZƗ�fK�v����_�x����x��. Zu��k1m�3�{;y�ر#3��n��,�r ����|ޞ����VotCc��w-���G½\< ��z/_ly�nk�x��ܗ�Z#..�!H=W��a�[8n�Ӿ����M��F���+��[��F-�&�cl���5��+� �u�#7P��1�	Gmq�pC1	�G6�
R�!�򙭼M�]��6�pV
��:kLb�,��1X��؊����X������	.�sط��u�2�3L�1�d���l��q3CB��ƺ��-�&���As�],�4	�45�e��d�f]����5��a�Ih`)A������~�:�=�g'�Qwu)��W�y��e�&ޥT�`�P�a�`�eQaH��rNks������a�[Qx��j�b��S!���:i�*]���a�β�KP�t3R�� '�/�V^�-yKp�fdelÎ�n5�����,}�O���}��^��*e	�2�I���(�-o��0�K�@�틺���~�������9�'%���~��T�S�313]W1����yX��$~@�o���G˥�����hfDZ�S(�#(��$:��7;���w�;�{�1y�̹5���y��ݞ��_?�O��haXU.�ё�c߹2�́�7}��_h]=ž�-��m|���֒� b�R �4�/�S�f����0�5�5[�ŵ�.�Z3�9�w)49�o}��f`s2����w�?������̬��K���݆�wGz;z����|l�5�.��o���y�"�:j�����Z*.V�-R6��7�Eu S��Z�C�hʗ���$�
ז+:��AY��f��^�ٮ����/o\9~��&� ����+8op3��a�y-�
���˲� +�19
~��Y7J�zr3�B�p!������y�X�1y�̽� ��%��Y��y��y�[[_L_W뜜�~d��۞~�5����1�q���uhV���O7��� B@��w�>����M���̣*�%�a�_mLtu#�\@PA�H%(�kgSw7<��� I��F��\_�"�c߾�p~���LPֲ��8�R�c�d�f�h��4i��	C�͕�V)�s��C�.԰�	F �6�?o���Ν+^�t�Y��*� ����_}o�O�0�f�.o���߼�}9���J��n�E��>�繿Fd��$�l0*��L]�[s�T����_y��y�?��:��50p��l�1��w1��Ҟ�[�z9u"B>��!��� ��G�Ս��h���=��M�dF-���R+�����9Ғok)X�B�F(X��@4z�?T����`t4vn�[ힾo��+>��N�9�AǂL�AIS��z��޹s��:"&"!L���N�/�|�rR�`o>�}裏�����u|���2`H���~��{��Z]�Wa����������u�9>�$WF���F�T\߾�����5��
�b��^@�:W �&�q��X�1+�V\���y(��9�B��:wԽ��M�:e�7ܟ���23�qr^g��$� ��d�S�g�bߑJ"T*baəWW91�_&�d!�;�ouF����uu��b�Iyr�v-�z4~��gy���LDK�������'0��l�@����|>]Q��-���X�S�))�������eɬd��V�վ;�"2.�"�q�~x�q�@�$B��B�\D�� M!t�F�d+�t�26.@�< �>t����+�6}��>�-ш���8�2�uh�/��գ��3����iL���j�2ݢ��/H���ڧB��tv��xfm���b�8��h�]�����S�&�>M�@$�|�ys�g�AG�	������l���e��z����=яu�T�ʾ����}/�;5c�ܭ�]p�&R[x6%��8��b�n�fh�M���ۥ�w�!=$����j�
PS3"��|Z�r妶�y�~d�r(t� &6�1������A	�		FHS�v�a�߀���<+c��V��Y�u���̹���*�7���B!D�LD�GNN�I�ޭw7<�s/�ߎ���َ����B�N�S
A�H��u|�Z����Ͻܾ���c�d����&�0N Mt����s�a�(��<�D�1&E�}yOs~�˙��GWY��M§-l��G���=���+=��=y�8��f�aDA�V��a{�-x
><�FFV�j�\L�nK�V���ۍ>�^N02�%����e�M�-f�2Ѽ@�F� �.+�JgI����˦[)������!��
�EוŖ�Ѣ��v-E��Fh�n�ii�Bй�p,?��g���\�������]��L��m���tIb��W��g���v���Q�-";7A�b�F��"ī6n�B�1��k�[f�b=U�e��.�]n�mF����UqMFZ�nZ�d�kMc2��~3�z���W����cp����=��˼�n���ϟe�:F���QQ�<����{�mE�p��ӝ�s"����?�t� E�&��B�D�4Z]Zg.(���Y�f��c��,&x$Aнs���Rf�(c���)�=��>}��s~>����W&  M�o�us���d�u���b\+�߻��O��ӓ��� ��q/����W[��|{�Lf���>�}�km�nK4X��w���:<ߺ��)�y�恐���Sѵ�#��"�2��h%ە��l�y�}�>���'�^��G>�;=Ssu��⺾M��(w@�-��z���O�0ÖݓU|���<��W\�:N$�g}\���c�]_�y�YW_r_�Ч���i�rL����.�e��4^uC#��Z�؛qr�rVal��=d�O3>1�
f!#3�c��G�}kcd��ٌ�K�$��y;<�[�br"P��D�2��t�o�h��dV $�- 2��IJ�ӟA�(��ɥ�+�|8��'j|��޸��9u�]��z%�����*FA��:z�G3�1���/L�O<��f�3ۈ��ϛ\���4�:h�Ӊ��N61!/r�����}^��n2os�77_Ne̻D�H~��߭��\�r�U��S�|{���|�f���	-~ߧ����������|w�.�+uxݜ��~��}�0�;�O�B��=��<���.C	>8���V��O��#萍z�����^�7��ֿ!	IN�����<��u������-h+��&"
�)D�唲��f�1��.�����i�4���m[y���~��70M��E�_ᄦ>�|��t�㕏�s�O���!o�3�ymmB�u9.�h���U���̣9��`���;���B�{{�|�Y�7/��@/�~��sￃk ��$����ޏ�tیn��#	j�7ύx�;Pq�O����N=�D�
"�{��&y�2.j<>�����=�t�X��Z�Z���;��N���	�3w��,I{��xn�?(�LL�Pǲ��v�~<(�pf�8g�儔=7�ⱎh%�01P��W��I��[v������&f�$�'�O*�fK��2����>޷���?w����3�U�e�"$=�����l��@����32�����WW�f\�d���s��y�/���7��NC���_䬌��gZ�c3����n7LZP,ٮ�V�3��L������%͊cK
ċ�^6�-���}����k�|��6Z��� �I����Y�O�Q`ǡ)hy�LľE�]e���R$ �>�ێ[7G�~�����d�D;3�ӰK�Dt�Q"L�&$�vs�cgg&\��!�g������t�S�]dž4̺��2�wR�/o|�'����tl��T�_�a�տ bN�b����G�0��ug�dC�//>�M�O��r�@���n��E/O/�9�Yt��خ~�N��c�Q3��r����E���۪[r�U3"�U.M����k�T#r�	�h��1Qk���{<���Ag}�N�C�������W�.��13̼d]��ȹ�\�@��u��N��uW�ʋ��&���.�E���l�r�J��nVbÃJа�ĺ(e��V3�������K�>c� ������OO�T���N���L6>��q)|O�￶/�������l�����2��gMO���W7�77�����O���}}���pF�h9~w���P�x����b�w�Sѵ��Qu~�1��
T����x���f�ћ�W_|�}����{��YE��76  �Y��[[�{��"^I�(x�Ǻ#3{�n� O��Lf�=��>��s~�D6j�0q(/
�]���|,��M�R(�C2��ӹ��w����5k�Ё���3�ʈ�M�%�`���2\��@�V�RLWE,T�cc���-���X���٬�Cd����Be���4H9GT6��2�[�p��%���]6��(L�Sk1���U�fn�0"S) �mn`�9Z��h�%�b�������Zʹ��� 2�m��off��-��ٽf���Z���̸u-��.�U !�j�k��Ix�F���b̴9u�͍�����wI��X�i��n�vez��/���������n�W�oކL0k���yyp����=�/me������iO�J�ءDiF4Y]�+�i3D��c��<�D\�b%Y�7�t���{��`ҙ�6_�<M7�����ӽ=��O���7X�.���Ɥ����L�D9312]_���/�.�0_m�����H��ou�S�9&�`d�uK���Ĵ��K�2mo���E��]�E�&niB6����OM�P�)u�@�t��"b��2�0���#}ϵ�ً�ȿ������G�]�O>�ͮN�I��QJ�fL���2���2\4:@	���6v���q�H��ouɕ���,1ݬ�ۙ��pnkYX�ULܩ�5�kK~�"XN n�޷c��I
3+�h��W7W�98�E�z9���7�߷�wW�ϓٞ!EK�*aJ� ����κ��L #9�C�]9#��7�Q�h������=$��:%4��M)	�}����>F��5���k�]=�v������%�g����[ɡ<ޮ2�]k��7�Ԇ62o�6n&j7u����b,����AN%���
7'�y��>�YFM�̗RI���uk��9Pĩ�yR@�'>����"�>��s̹�H@2�}�;]�Y�7x
a�˸4Dʷ�o	.q� c=[�V���~���W��̬`;�����?@�P��)R�o��<|���|$r@�D�/���Ӿ��跿[��|ߺ�r>�I唻�J�)�5� %ˆؘ���h��k,qc�]At6.�(d>� I>p�������HID�T��}�ˍ��,9���(乱 �!o�x��}���]Z�R�E�[�����>}�>��HV�z7�����*�d�̗&·�q�छD��&�)5����=�>\���r��0G����mݾ2�5hć���S���v9O-�7��it�sk��-�ɝ]��e���[IOj�״�n_:1�\�	௠��˸�מ�J�W��5V)�c��[QQ��uv󜾷�s�N�u3J�s&s���#w2�2*��V�\kn�$k�O�7s��ݞ{�v�LT��t�i
C�Q4�!qC��Z1q�s�����g�G���y�VAj��35���.'����V��^K��S�?,�w�r�R��'y�|!s�#"�#&���s)@w�&쉱�^]�:���f!x}G;};&�mI�	��bt�W�qn��+Yq�7�I�Nr)�C���O���9u��7bL+������qg�d��M�5�1;����d�en���<�Sϸ�EgC�
ܻz�ۦ��[⭙n�N����?��.�n�?y'W!�۸�p�*����^���o8}�_�O����O͸�<{�7��׭��fN9��7T�j���o�l��zP�>(7�b$�1��A�yc艒k����^J���uܶ�3*[ݾS	=[���hbzf�a�='�3<n=��dwq9�X�+9wù@9�±��>���tY���㜫�w�=�E=ίn��ٴ��S��}�:��.ߧ�X�ҥ}T!�4c8��Ds��خ�7����N��S�w����n@B�$�ܪP�u(t3�O=�.:�h}��^R�;E��.Q�5��o���iVn�k�`lD�nT9,,¬���:���T�S���O'Uu�n��:�������T�s�o�{]��|��׆ջb�����/e{�{���|�x���'E�< i�������Ҵ�?XqT<������zvR ��bPFU_P�=��z�{����M���e��b�.��d��16����H�,��Ѹ�q�׈��'��7���������m�EZ4�{��ns�LW�N�+�b��ŸV.꟝�������	}���6��zyh�$�i��U��"=e�x��/��L�:����k�pso�� �Zt�6�k�l؃�?dyI������y5�ϕ����2��,��������*�y��C�b���f�ur�	���k���k���^�o=��sGf��y{QO�����l�������-�����Gސ{�cU9�V���[�'}�zK�yI��ӻ��+�F<���@�e�v��9�����F�d��w�-lZ��U��֕���]������D��qu7��A;�ՏgO-!f�2zYx�v�	��XQ� CY�,Nb�ɻ��@��<5ynE�<>�`>k_�/�Y�M8�_�(���{���L'��pc����?u���і�u��Z����2l�:�G��
���s�°@����cѸ�����3�ܠ���c(�;���R��Sv(=vA�=�n�+��g���邐Q���D� ]�-�Zm����OK��8�f�B-�<��V>�H�/zy�;�C�Ϻ䴊�����^�=��ڻ=�:ײ֧�t�U�{S���W� ���Һ���������
#��!<�2�/�\�l ����vN��s�YFM�2�L �C��w-��͡?��@(����E��VN=�2nJ�@��tk�cxʿ}1���w�$��`zlb�o�V�gK�V�)�e�4s�[u��&��BXݫ*p���������d��R��SLO�����x{�}1�-| ���^�g>�+F�N-�s�/CKT�����/ug�M�+`�|���s���a�~��T�3'\�����DG
	�	�Rx��[Y�/�����r9�r��%���|��w֝l��4L̅@��S&=�7&P%�w��ճ��q~0���_)��PD�O��{ԋ�Zz��DkλyJf��:�t�1k�G��lw2�Xڛ�U� 3G���яc�w��$jB����~|f8�����5p�����v 㒂x6٬�x&P�Q��/��v Ϟ9U	����0
��󾳰�(o�
%(�*eJ�;:��Ǻ�nrCz��ѴwV�d]c�a�oӞ�<��oXmB��#n�)����1�ˍ6���]���1x�uq+�Z��r�N���
QJD3=P�~[;q��8�i�~e��F ���ލ����3�𩤇S;ľU�fN>rK�L��F���1�[D6�o�� ��WO��S((1I�3'N���M��s��\�r����r3x��;��1�V>ǡ��11�|��h������������/'#�����Y�����~�ǈ�x]#�&H�^��E�>=�$����������;����6ЉYɊ���4E�d�-	���&!%�Մx���u�O4R�@�< �NҗXm�A�>`����_w������)G�l�Dc�Y�ve�BX�m�k����3Մ%ѷ.����A���!4����CAĎ�4���{�&�J�D���C��z��̰�K�f�`�%i;�em6qnԅ%�+�V��-��`�գ*L86o`-�X�X�]ʲ�.oVA��o!.6������.G�5�@�e�6�6-,��0�M5iC��d��1��6@/��x��7_-�:J�=¬7�&V�v����#�aA,P�Y�pܪ	*�j��^�%��s��(�Cf��{�?Zm�ǝ	���j�p4�@��i)q��ܻ\Gx5��'+DR�tԪM���d�z{�[�A�D)��K�.6�Ա���������������G��w�V�j�#�d|߻��9��l$ �s��峵��⺿E��_$���8���F���8�*a;�2�2��%�z..~y�2�%��aX�'�_V���6��)�ܙS�K�_2\�^�ݛ=���\�G�<�7뼟NU�74��`@�ٳ�y&�.A//(y�"�/Td_�3rR������پ�T��}1����̕.\��}Mm�/1�WK�ck4`��˴V�Ln7`�Kf�.,cY�����JTVkK�c��{�z�-�a�1���<���ᗆg�ܙ����F�³�����a�I7Ϡ�����PD�A3�ypLGXFK adV�{k2|����ş#�*���TQ�}7�a�4<bi�=9{�Q
B=�^�r}i�^�On�=;�Vm'ku���u�M�4�����ޢb�{ BLҫ�d�9�*�շ�f�|����n�Ў�Q��vv������>';_����*R���2���g�8�i�p��� 2�s�[�l�g�nn�##�<;��^"IA2����� `H���GF�z+&������5��>�:����"̓�<��JʿC�ⷿs&�с�?_�Ӵww�.n��{��5�N'�2Y��`F�%K�e��ܴ��G�f��^ƴ�5l�J.��w�~F�yV|�-��Qq��َ鷿�bȺ/drM���t$ﾎ��}��Ǟ�
'�x�y������|�h�$ �]>�>��߫'��|�K���`�r����"Lğ��'�a��:�6��en5�c��� J�i;V�LFj�5��5�#��:'���5��~13�wI�<��_a]x{L�n�CPwP97�q���ݲ�6yz>�!v{����\�Ϛ������W�1W��z:F̫�B~���J}�2:�;�v6p:$�]
��y��{��3/��7��յ���]_��1d_$˛�� d]Z�>]_�b
�)(��L��K[z����s.��3-���k�F�Td_�"�m�y)!�{�OT��3L���e5�`�J؛���k[v����Ō�[cp���I�i�n��nuQ ğL�*&er�j{��k%���Ա�2�Bdm��t�vvo�=C���f]�&!<L�\]G�8�ɺ�wH,gW����WVN��kl�6���@ ���H�S_�x�Xl���^����{b��J���}S�~�쨸�|��Rʋ�R�����$!��?�}������=�u���[����Ѹo�	�l�$2��̟a�xZO�G��1�ɴ*�*��c]����|���F��KVvA��7�w^�D�
$�Ho �����3�K��Shjx7!����b���9�e����G���۟OD~����$ ��mr���O=<�O��Ԝ���Q���[�[_x	��H߇;:X�J��8�k�PNպ\��.�a�%��]d;��D��u��,�w��*HO'F�Ⱥɋŏu����$� @�s}�Fl���}d�DrB�&%��DK�\��d�&\�e;��ꎍ��7���ӓ�972�@�!����*fe1 �3"f$uu|��l���M}����dz����w�o}Q����	���U#��Ĩ��̿+����Ξ�:3�7Y1�^Fs7Xˆwv����6v��I�I

��!0D�N���;x�m���~���xɿ|�xe^z��+��w��r/���ݹ�*.ɪr �Bh#�[:qV��P����<c�p�gMGN�����������tk@�ې����Q�.�f,�r�2.�$kd�GJY�v��"�+4փ2!�(�.V9�̌�i3-�l�m&e����&׍]����R3�b���TJ\�h�-Q
[�R�ѥ+��]��I��f�0T]�J�LV�����0�Am��bi�uK�1(1qw��2��i�c	S!`qZ�m�2mW=�m���t����j]y���/ �,+2���}޹�	�����ُef�1���7t3�x  1���y��ϖv����B�x!�-ԘLI݂J��H�Q�ă6p�K��sl��Im]u��.tu��]^/)��'8C�mԽ]��j�k«��=��v��K��N������G���Q�������e��)�T�:߷���.K�����t�Q���ɺɋ�y�,��g��p��(%(�g�f67ޛ����fd�nk��|3! �ތ����t�����x�(�!�I�2�9�83,��][��|��9踾L��������&�\�D��<<Bw�2&��zqees7&��:�����3�d7e:q6���Z��JB�$D�(��:;�4
5��Ћ�F�6a̬�a!���i�Vrs�;��ubÁ�D< �>�_���b�۽=��� >�H�y����Z�`,$�&A���L��Í�S���[^���G��N@�y��Ǒ:l�σ}]��g�C�H �^c�Ub� 
>�>��#S�Ӕ/��|�
VG���Sd�L�p|n�%ACJ�r��c�/֘�T]��Hj�m_���.��v�]Mf��t7�@�0N�_G���N[���i��B>��jk9�N�_L6uó��oܟs�����|�ϋ�aQ�kL��f>��Ǜ���'��r�]�mu��c>�8n�Œ�U�#&'�bS�����{����l�noޛ����M�� N?u��}~w�����6�g�X��9QqyE��rP&�d{x���T�,�߇��)n��x\������DD",����]�XbjjI�H��XC�Vl4#W3hX�5�@N� ����YuE�K\޸�E_<-�tV�-<M���E4�|^}[irL널 @��2r�0]]Q?	����ׯ5�D����u���"�'f)02<V�j���qb���+	0^��7��&G �0*�u��R���ng^���|�z�4�J���XI�⑰c{.�sdS'�G�NLԯ���k��^���2�@M =DI����lXF�=p�3� ���v;���L�1
���@�h��X=C]3uD'L��\R�7�Ǻ��i��g�c���^K�����b�F��� �O�A��4͐���U�פ���xw������X&���ڞ�̝7B�}S����/��+ݳZ@��9��Z(�Ù|遷s��_8�S�^���6��ԭs�^	�;+��g^��_�I;-�{��x�
�<OOqK5��u�\�4Y����~IB����Ui��iu匪���tR$���0n�س#�N���'3��%��ŋ����|bǝ{�*�O��ͫ�Zx҅9��ɏ$&	i�E#��=q��U���������x��jwJ[���m�I�8�O]\֞4U����ZH���V��`�}0���D��q���Xx��^�}Zx�|<��$� M��<s��p�҉��T�^M,X��Nl/K�!DBxx���$Ù�1�L�W���\xX|M�x����;sKOw��)�AS�8DT�j�<���}�a�@O��������DxI�@�B3R��X���y`0@giZ�W̥�[1/��K�X�}���j~=���J�1�@��~0���7{��EU��a��7s��"�\")��8��bo�5��/��)8BF��:yN��+Ou�3�Z�E��L) g}�
����)���Fb�{:k�Ƌ�����Kt�F�U&�"v;r*J̄t�SB���4wcLi�4*�o��z�{��zX`R�1 �LW6���s��<l�]]1ZI��y�ҹ1I 2��w>�bȭ"�+�ޕ�3��!���X�=Z�9�t�L����}�*��p�:�L�����P�� �9:>?���}�?��J�b[���4_�V���n�ޚ�{�4�m>:�����q�7�^}߼F���5F].��zvO~�܄I�oO\V�|�x���)i�O
���+Os$5�$Yܫ���g�}3�be��PL�֊L(���K5���fB�00 o���(�}����+H���U���p��������e
�v'&�ϯ}*�r6��or�gz�^"���SЈ�ќ�+���&�U���_Ƣ����sv��{q��v�b�]}(Jr'v/0�/=�z�x�\݃����q|�n�k�Ō�Y�5m�0���c�yf��͸��[���c=��k:Fd�y6wH3T:`��]�̂�]�TGF�l����ytR�j.�fso��l`�q�NN��}Z��ԋ��뤫�9���Vs��	�sg�c��.
�2����yf�Sa�W'��[��z��j���ɮЦw�F�}�a�#�>મ����s�(�閎k��	3ˑ�$E����
ȗ���rzo��ƺ�᦯#^��rE�k�U
"0�j����\���.�C�������ވ�{�T�xL��?�)��)�9�$A�,I�V�{n����u�x`�/�7���=�<�v�8��{+���M�:mQ)�F++{e$O�UV9fF�{X�қ
���Ȳx|~G���oay�X�N�[k�i����,D���Y��t�m[�0�.�&[�qc��{o��v�ϟ�8���)��Fҫ��]RV[���扜'/��Dd�[9���]*7�K��ڌ�����w�����m�`�qq�:{���k�\����>�aϧi�Cok��t�ߘ�;gp�|�svgS�5,�Y��`���)�{~��W���c�ZY��������f6������l�dd)�{i�k������.��3�/�sT�3�r�@���9W5]�6�0Utu<NE+\�
y7¸Iܬ�8�ɡP0<��޽��|*8�3�����ޞL9Y���+�����8��M�뽞�����Ͽ�w=q-� �@��V;cfZ�����
]X�-��&s1	�a!��<����6�p�J�Tl�%����k�v�KC��1v�����:.HCmY{h��X�v��˙@ј@���#jԲ�Y�ʷ�1�cf�7F޽�Wp^F�V�8Xfc;e���s.�M�v�=u˕�au5�fe��� X�B:� ��.�[���f��k p��^@*0�n#32et��mW/jS\6�m���G.xv-Nb�Q��n�iIb6
��]���u`vH���X卪6A4����k���(P�R�bƆ畷C������l^fׂ5��h1#�I�֔(��mcn`�d���U ivf�Q
W,��@�]J:����tv�W,tf%�����n������7�4�ٴ��e M�]��1VT�1�\)���:���j�;JX�LlQ;حJ%�(R�s.֨9�Z����6�8�T.`�L��R�a�3X�l
6��K3u����m�,��RkMS+�b6T�-5tD�!EĲ��Guҳ7�V��7�� �G9.�ǴfUQ�]�ա��)d(�lYvI�M��76&�(q�k,,�q
�i�*jۣ/���XDF�0Eұr�1ƽs-���1���Gf��#��"\�%B��V6Ԙ��pu83��T�۰���6���Q`9�tz��71Ku
���V��"Fj���b]f]� ����1��Ι���.l��V]�m�g��"�l�Jh݂P�A����n�r�L.v]Z��H]5�-t�ZZ�8�`�	���[M��B]u��s`U�<P&s��8ڳ$�l�Rjb�@N��jM#�`�К����n9&B�١�
��Ŭ)hc5LSA�ve��n9��fFa���-ܷ�͖�q�ڔ�nH�ƚVz��Z�R����uI��cz��S�����W\��c6e�.�4�H�3�Ik�lݘL���&�At�g���B�4��H%jF"A�d8�s��m�Ě2��V�\R;�.��%�-%����=�I�\q�u�S̠{�G�w��U��)i�_y����M3�iv�ֵ�=ƫ�J.�x����.f��Jl��w�SY:�f�������$��T�-|�3��;eK"JoU��uXƷ/L���܎j�g��V���K�zŔ������
�Gj�/%aC�������ݴP��%�kc/v��]h3J�#�45�>�����,�;&�\�ǽ{���$�)=:Ԉ ���H��f�ֶ��b��A������D�l
�����2�o4=N�Yq����~Ǒ-�z3V�
�f�������p��Zkh���;"�tM8��㡡���+�~�_
<|���ּ堡����YU�Gۅ�t�D��3����q����yM��O�W1��K���|���T��p���
����׾��)[_��==xي[*�fl\̣V�Z�utb�z��t�c��'`�����<���ŪF��εz�����3���̉�^znwj�� ���
}quW�M����̭4��-�����+�.V6[�qr�)���k�o���ui�O��Gn�%�Ɏ�=�=R�8
K��+#���&����lc��OV�p��0k��s��Z��Ua�b�8�6�8j5��A�wkXA�Ǵ5��KrTT������u{�e"���M-z6l�=��,���A��+R�w�	�[�B`C�t�	���qe�hJ�e����j��\:%%�)G35Ë�K�1ʶ먆����m���`�hM�k�D,R�f����b�U��yHpZ�k�W	O��z���.-���Z�q[Ҹw6�.�&��I\s�]Z�\����n[a�b�J.������Mm�ל]�f1e (�@�e�[mX�%kv4��:�f�`D]e��ke"��a����])�B*�iXE,��<��|���C�����\}晛����z<�/_U��6ލ�����_r�\&��s���_v��yY��#�q<x`5���x��j���u��2ٕ��]4�����$�`��t��s����I��GJ��N�f=:#i��S4Yv)�6Gr��o�~�$ ���<uOqK����LP�t!K�#��/XI���s�-U�&��9�Y��Z(�����KJ4�=�"��a7�``_(6;�V��30'R<ʮ$[���Eh���T�^NmӀ������ZQ���[��V�OO���N�ቝ-�s��w|�r���yR�(O;�=a&��5�2[���."}�M|/P����D<D�&d���i�'~+
0U�3Bo��33�{���� _Ooz+4�|nN�KJ4�rn��<:�OLC���;J��1�2�U�Ѹ�u��1\[�6Z��L�5���Ӝ�z;�w�z�Q��n��;+�ߊ�E�����֊L(��ҿ$�V@������zkJ4_|���jx�!�w�Z�b��i�zkeм��c��E�>A^}u�N!g
 QZ��'��R�-Oe�>P�<�Y������>q�m����b����TQ˛:#E�H��M��nwoX�wznJ���H֤��n�������9�vLU����[��"v0S�T�ОE��_x�e���T��J�n�XI��u;���b�M�+s��T��x%�<��LL�b��Z��^M,[聆���h���{:"��a��ձX/K�����L�DÒ�]�<L�-(�L��0�e𳧾��<h�o�V�-����~��I�$�R39�g����qb��a�;<��P�3�/|��ߞ����:ed����^������KH4�<��a&�ܓ���5իv�5h7Q��e�-(f�&�a�y�ˋ�H�V3j�������N�)�C���C���H���J�<.糶k��(��l��y4�U�s$� ��KO!�]�*��l�hvP�Q"R�"D�֋�|<lf�Ky�vN$������Zx�|<�qZH�_�c����s0�� p z~>����oĶlT��3���qb�߽�/|��ߞ��|�~��vCN��(�鉈{�ҜM��ސ��D��e�Qc*�%����E��7d@�wQ�[�3�P���>��M�e�"=1�z=ň�ǽV~�����F�]��]����*����!{M�R��A��(�>��"�i���
`�:���=I��I2�XI�&-���=��\x[�eeW*�Q��T��-ףNd�]�������^�:='_�{�>�:�t�s*�ZH��{��V���x�V����g�ǎ(Y��QXx�|<�iZH�_�l��~��Ca��w&�$eĮI�����,�┋���˚kS:��4'>9)�S����ɪ����cӣ޾���=?}�zk
0^��7��!�Xf�����^�������u��e"�ĹgS��'�݇����d�h��ur�<.粲kU`����w�,���Ih	a��7��RD\A4�l����.�;��ZP���߽5���(K� K����J_qB��z^�����:���$�"b];ĕ��w�C3h����Q=9ʖ�ɥ�k~��a���9�Lmʾuj��.�}Ei�מO�����Ñ>4�H��>	*�2�ߪ�a3�D��^G\3��Ȇ'x����#e�{qonU![��U�f�һެ�	�'s�K�������=y��nOw9�z�|�Ufzɧ9�f�B�{���d3��
=�2�I�&aL�2.�>6=�R�(�a�*���J4_]�+Ou쬚�X*0��˹R���.<�T#�:�A��j�ym�.�24K5��� ��n�b?$�^�����[�j%�Ҏ}??O���Y��V�`������O���z�C)A¯�K�����P�5���C�H:�/Zx�|<�iZs	��e�w>�<W
M<ONj���ib�oޚÒ@�}��c�}�	䐒f&+������^���[9���rL(3 �(��"��E�}��Zx[�񰻾��s�r+:�}.'����3����H��ɮ4Yj(�ʸ�y�I8��1o����
|�|Sl�x�א�0���
eP�G�����h�3���(��+�s�t���A����f��X������r�g�.�#�ϼ��(�R��Yz�R�ΆG,�I@@����2Hɛ]5ր�hS��S�e�Z2���!H]�R�
�Ք���2�.73GK�攁5�ʐ�YnI��X��K�:c��zzs��]5x��c����^`J�2�Й��l�Ye���L�I.�^�l��an�M5�X�$+���`Ie-.�m��Y������򅆎j��E�b��v������mw1�Hf6#142�SQV����*KPĆ�b6/�?���k5��܎��d���\����N�<6��y��D��ik��@_���cy������\�Y�,���+�k�QGZ��B�at`�e�eѳL^v6׳�V�\�gz�_[�>ff&i�,����q�8���j������sU~f.$��N�x�ҍ��q�fJ�	��ZxY�ⲫUā� dY�=sK��8�g~��L�z�͈�97	ӯ�'C3��5t����HI�4j|3a�Q;����A�>�Z�����;3��D�緊���gӯI��z}ޤ3k��8ٝO}�̝p����I�q?��5�/������������s$2o�k>�o*_q�8�����G��1�/�������s3�m��ʸ^4�ڞ饺�ib����J0_y�����u��C�[7!-F͂Rʑ)sL¬1i��npsi�l�Tv���8@�,��[�snM���Da�����2.�8k]r�Ə!����&G�����H�]ʸ�w?è�v���c��zLxt{����{��9cx�a��]�q�o۵O�3@�r��[�U>��E���덻�����7����n�	�^�$�9����s���d��
���x���,�:q�3��4���|�oh�~�2���
nk��*�)�R���Xjk�p�&���>8���@�8t�ެ��E�X���W#��-S#�x�������

�2�AR�LLʥ�P��|�XQ����j�<rL2�$	w=�W�Mp�i�u;�-����S{���*F��^�:<>�s�N�=��*������i�T��Z��4x�D���Ѿ�+J4_<���N<J�H;̪�E��}�Z(0��!H��B�߹R�z8��_MaF
�{�o�ZvOO��������74�5��V.��h�Њ������Ι�*�6�l�Fau5����{�7�O��2�w�z�W�O��o*ZA�	�7�z��ߊ�7��;����'g����~���uU��u=���*�ߊ�L���4W����ǅ���Mh�O��^o������%�T��'��OOI���d�p�+�*҅��3�y��L���K�pX/v 6>���|����"ḏ{��;�UuC%�=�#ƴ�{�D�s3�'�|4Z{2����ox�WCU#T�������'� W�� �V��5z���f��ݞEz�lf�^y�� kʲ��qy���Ƞw~���i�[;�C�Q�dOv\S4Y��%�����DL��b��o&N�2�Y�����|t{���P�k6
�L9$/������N�;'�^���Y���v��"�/^����sJ[�񥜗;$=u�q&��z��ZP�����V
i���n�����-Z��,���@ 0R�K�.���A�6�2iK�3``�����s'V�4�V�F�z^(��o{�3ZQ��{�Ҵ�f���Y��03�O]]4��N,Sc��������=�m�iɐˆbs�w_��^����?lR�(O��a����!/(;ͬ��%J	���_#�V{��k���S�4�^Nd2K��}o\Q����{b+I'���iײ�m���-����:o�Iy������ޗ�|-�o�k
0_u���ܾ��2��ө���D�]��7������
�m��5<Q���e#5J�㒟u��v�tgC��٣7���o�N5!�Uv8mkVY�V�h��V�P`��m�� �,����n�֨���̻�
��A>4����cӣ�x�]��c(٭�Y��ڞ�����(�{�d�/����ʊ�����zk�>���- ̛҅[� 9B��Q� �
-�����Vé�U��Sf�F4��]�%��f�O�'g��ys1�-�����'��������3�Z�����+�2�@����<)���\I���ƺ��x�
]I2LV�-(ܝ�kd/�}��gٽ祅|,��XQ��{��ZrBJ�I:�|+�z�Aᚪ,�J+��ǧG�}ׯS�jz~#������K�`e��|��=q�a�}�yO�M>{�㡤[E��-Jng��$�	  e�N�t=i&�����i�n��߫�X/rHe $	Y�����G��{��jj�k�p�^��=����OOs$��kE�}<Voy�iF�+7���/�K��(���8�})����(�dh�p�'H$v>�׮����$
�j�	&�^>��\�/��d����<`� .6M�Xl�j�&���S	�T$&�45��7�V��nBhL��0��f�.��Hh�ݠ�a5,-�Y\��)UZL`ו�%n1)�!0M��B1��Rڶɴ�����1�A�3IIubki�\���K6v�P�%�k�"��`˔�V��]mC �#(� ��qJ�u�Y����R��\-l��kDV�#��!��SmY�>���G�G��
�7�)ɕHo������)��q�'�G/B�#�پ�xh��r����-�xn�5:�}�}?�����M��."5Y��m�i��n8��I65�m5�sk�\�X�Oa9 �;�]N�i2��vw_����Ǭ��޽"xvy[[4�^M,U���&��x�]�{{���zt�u�Os��.w^��x͟�io2N��	4�xO��Ei&���o�i�n���V��s3	&����狁� ���4���,[�領�<nm�֔s%Β�>;g��z_O{��g����!o���Y,"SM��9$X��o*���!VW*�I�����Y�&��.�?���ҍ�=�(/� B�"&eDJ�0G+�dW4�x�±%����(O��Ea&���U��|��x�d�0�)�!�!E�h5׎��V��sGZ�XەK�V���k0S�� I:���ֹ�Y���|N�?T�!��!�̚�DM �� O
�_Ep�ϧ��u�$�ʈ�f^��i�+6J�KM4���y��՞���d�L5�wwI�T"A #�q��w	�4��i孝�Z�XЦ�p��Tl�W�4�K�'M�w/N��p{��`ME\�Qݞ�g���6��[D^v���y���U��? 8H<l�)��V�!���&�k��
2��if�3!2���'뿁
l�N4�)&���m=���|4g��f��X/{�(I/�ZY�9�K�(O՝a&��k뻸��//	�DDIZxY��Be��a�W����WE,��6~�+Ord2�`��x���WP���J3(Dʙ*f+��L٭}j��i�ɐ�-�o*�9�V,<n���h�I��7Ý��uNS�Bx��-XV��e�Qر��;��)��.�H�f�^�]$�8����c�f5h��������j�(�|<���,<n�}�0�Dc�����t����iB�@�����w�2V`�����Nfa$��3�ܫ��O���T��
��b��J_O㿢Y}��mU�_	<?���.)�E�3��Pf�����p���[�|!F��KQ2P���3sv�s��TS}�8��}�Z��I�|���n��[����:<��}��o�f�dUN�OH5��,vrLc�v<#�r�A*��7�6H�;�S
�ȃv�}�C�3z��A�͈�tsK��H�ub�T`T�wK~�V��Ik��#�������Ѻ��F�Nh��F�O'=rr��oC��n��}&��0�g�U\���'�quM��Q�9n�r�nڮ�f9=R7`�V�yN�u�R���ܝ|2p�["`v�ŭ����{�~���4v�������d�(�s�����3q��-��瓄�ۛ�V�~=v��l���/���eI�����=�`H�C]�m���0�_v���T���|�1�J�Ǳî��}|h������z_�C�iTq���<�M+�k��}w�ǫ=^��r�1978ۙ��&���ri��z�VL��?M�GɁ�o�Ԭ�g����澳$ܨ�T`�S�9��ͷ��ɥ��ө�w*r�X�7U��ܘ!u���,�va�YWF�K�[n�p�6$�V�.��]S��gI���gQ�N��6sb�o'����U��YlnA�r1]��Xﶜ�����֦����ȘG���W�7�����ݛ潯�sP:2Y��4��\�=������=�1��+��i��igl4�� 	\���#��+�Z֑�M�����mM�_/�)�#���\}e�p��>�=��3����6\�M���{�*\�c1���Ƚ�k�G嵤������|�T�Eo��eT냲���oi�ϭ��ȅ v��W�Y9��-�TRHt�+BV�TqK�l	�t�G��[ѿ�����}��,�?D�E�������+>����UQ�䍋�߼K=���3so���nwz_K�{%�+ղ���{���v�f�B���j�^��JzT�5�s@�R�qw=��9�`���TxcUS�vOY|��g�{{�����UѾ�x��k�3l���K;v[����F�L�r%݋t�Θ�����{�bԍإ}�\#�QM٫r4r�sf��w7]����A�5�Ԡ��6����p��X�YK$�h\9x"�.m��I�7a��+bE{|���*$��r�ߩ����d*�3u��[��Tu	ܐH�7�(ٶ�{����G���`�~�@=�N�޻w���]����ا���Uh�0 �j+����-Ʒ[aV^������7��EI?]`䃼��tƺ�Ki��"��|yh���:ׇ��"�Y']��9|�������n��˖Nv�>�v��s���i�LN��v�K���^,\l
��A5�̓"���j�CZj;�L��j��5�1��W�|���]x��.yo��v���Ci�D5z"�Ċs ��3(��m@og�:nv� ,�]xI����˰{m�	�+^�C���q�4���Y}V�+<;��t'{W��c�������o	�S�NM�3�x��#�i�7�����1e�!@wZ�sع�0�N��Qb˟Ln�4��17��lB����w�+^k.��=~��=��7S>�I�}�sH� fN@�9~+	4��μ�u��ó��w{Zh8���EUh��d�4&��ii�
o�UaF��sJ��Ó!2N&��~����=�[�e�b�F.gS���V`��'h�K#����ҋ�W*�x���o�XI��ɡos�;�"��
�.��.�n�ɪZ)�X�@^��͜i��Cv�q���$��=��jQ�:gV��kO/}\�����X*0�y��W&C�� Lx][\�I0^.:�Son��ں�;�����{�ק�	��OZA����zk/���+L3k�'>7�ʇ���S.<K�ƞ3��4��
���0��2c]9�=ei�iE�����F�#TDQ�)�gS�<����'��� �|�޴�ED�w�XP���߽���{�f�5tTH�"H�C�S^D2(JۚEP���ICIt����ْ��x_�t��"D���	S�>ƽ����r ��a[6��稍������ͼn���lq��D�Mz�G��b�<�^�\8�I[Ÿ�!N"�o��K�3 �/�A�=�}1��fD
i"bW��E㣽�X@���:f�]K��^Q;��K0�W[Z�/�L���8�f����x՗E�V�\�+��GM�!vIcE�gء��;��z��`�M
+*��p��e�dQf�E>����q\�)BL��7��<-(ꑝ��
"!)(IQ34Ȳ���h?��Hx�1�t֔h�L_l��ݯ��\�j�$�Ɵ��#�/D��*`�ʡ��#�u�Ȳ���f�$��d	ic�^�+�&��[������˽eڐf7J�u������eeo{���i����xج�KH0�J\BK���+I4^:)�DK��
f"b���u���^0��HiC2�oܩi&���������+J?'��"p�8�"i�^�]����,b������*���i���f`h�u)��yֲ�Tt�u��l��S�w*��m5h1��n���#��TF�v.ѳ8��k�m%)
�����h��.�PԹ�Y]Ț2�5aMe��Ct�Za^��^�*�M�:�_^��4��:�҈��@�Ϊޙ%fm��j�WSTe�%7BVh[v�BLF����с4�6Yk�].�F�]�m#@ɝ.�%%�K4˭�m0�[t�{G�1�[J%�J+*u��9m�LlRǕ/�~����yU�x��*�E��2�Ei�B����Px�&XkdbB2T�1zL�W��m���~vzb�矽4�u�<����E0�� �K2ZJ�a�6�bƎ����<�M�v����{�1�b+�f�"
���(�:�h��u>�\d�x|��+����I:4�ZY�+�EX��E6>�d�!!D�DL�f8Cw�5��\2i�,+��=i�a�ٿy�F3g�4��d2N$������:	$�a�T����/��Ea�a�u;��^�N�fKK+��R�M>F{����c�^���.�Eg^��ϧ/)�s��߫��^4���祥|'��U�rd2^C �ߺk��&�Gz&a�%�S�(��y��Q���K0���D�_��+O/�ޮ�������v}$��}.��^Z������g�j�\�l٭%������))kiL-���NRr�$	/]�ܣ��Vܳ�ُN��_}���L��V�a�a�u���0�C1Μ���ފZI�����9L����<� x��(�P�[�V�۶}qԴ�U��}��[�ћ^=o,B�(�=q9Rl3P��|xe��$z�C���,��Bf3���ye���;V�-3�i�K���*���y7�;,�Η<��#*���ʫno�z���Ν�W�S���Uޕ�{�B4f-��"�3yZ�����Y���HKF���

�����r«עON���~�&0�+kf�ra�@!��~��֞4_�����)�a�DK<�<L�h��I��%�=����'���i
��V�i�a̐�6��*�x��_�B�CD9V��x'�d�ǿZ���̝�d��q�i����x��Җa𹒬n^����%��K�IK�r�5��.RSl@��T�]"M��@��t���D<���P�0
&eW�����aB��l�l֊(��د��+2ҍ0������0���*�C���R�U3����~����0%���_E+ ҅���V�`�^O�+L�ec5�K�_�KZ�F��[�����������K8GwVE3G콁�^�|�G���l�xW��� �{j������wpr*|���k�����f'�%,$����ҭ�>�mn��J��o9���Ǳ���<��S���a>��_?r���x,�͠%����|;�n5P5/졙H���"��Y�r}�X/x���Mo�j�\��zvy��zyH�ѿr�$�x���k	>���E�I@	�ݼl��4��O�6�-".a�33L�da���L���^ }�=h���WW=, �����+
0TsO�>�e.�o�F���올[H���YX��\Y��&�cZ��e�a���B ��찮y��y\�f+OO���U�����^�aB̟l�&Bf��E�;��������B�8��gu�:<?��;�R�L��e�յʸ�E��=���aE����E̘o��4��;��wpft���^��=?�_<������Y�z��3!j d���=h�i���vu<;<;%O��{4Kxl�1���:H0f������s��Z/|nz�RҌ9�k�q�ܐ�}�B���{�{ܖu�У��z�\J]}ڈ��@GnĎ9$3�qG�M�z���߼�����.� �th'ޏ���k5��ܞ�����O:ʎ��I^�\mĺjϵ7]�8n�����#c�b��Ȣ�W�B1Б�&����$Xx�߽5��I�03{7�z^(��v��V�`�=�iXP��ɺg���
kq	��Wp��ItN˶4��\,�RRR'uM	r�����1���j
%K�(��Q;��K0�O9����/�[̐�e�
3��=h�i���u��A�.L�3�����=��{՜�;xd�Ɗ߻�ZxZ|]NqX/|\o�Rә#`b�O��u%�10���/\Q��򳢰�a�6w��$�M��}��K�Ɵ
��ʴ��_��]}�3.g^	<�Ig'����x�Q�;���L(O����reN�|{}��
ϋ���	�b\�	iy���<^�|R��9������ �Q�=�Z@����l֋�̵�7�G$>�z2vg�����.�<%���w"�>�<JK�$�\%�qz��.�3������P}J"�Iwiu+��Z��؛hz�{=�ZM�@�q�50��W9uy�L:�X�f���!D�Vh[���;�&h�xm`���0���]#������ں��Gc�٥�m�T�p���*bk@8�iB)Ж�4��eŉ�FR�v��S��&7h6X�[R6u&\$FXɜ�f���mj�4p��[H�6��))m�`��I,��U����DFؔ&���*J���8�KolDY0i�L=��5�uNK&�>�gI�M`�;�."qlh;B�݂B;�=���_��`LF�Mf�k�L����]�fu
�`�j�M��v�����'��|�ٕ3�
�40��d7u�L�daN�Eq"���3�f�Q���\���O���0��_��RDD!
d_��e:�3�Mn�|-,~:�z�A��XQ���y�i̐�X�^4V}���ǁ<�$J�fb%W��g��j�Y��u>9�(����(�x��tV�|��L̛[�U�,��vy���VUv��|.���ZQ���[�aÓ!$�@��oWEp�����2LS0��3*�4Y�7��W,���̎߹V�-(�U�V�(��lR���9���S����*� �L�RJ�s�M������6ð��96�n5�6i~t�=��4ID�HK�5�/[\�������Z)0�{��\�2�0 ���wz�+H4^9g����OD�D�a�a��{�q�ۈb�0��8���B�t�^���	 '�W����>�2����Z�>�{EfD����Ӱ8� f!W&m������TLר}�`}���+ؽ�t>`g4���=�a�v睌t��M��� өkz�?zQ��~�ř�T��O����֔`����+Hm&�	ώ��P��A/#����I���W=,(��^�|V�90�O�d�q�~�ZH����٭x�}�7��jd6^��<�Ig'�$�<�zkI4^&���J�z�xÓ�	Y�w��� ��N��L�(�S$��a
��V�a�a�2�f�$ ���U�x��;�����d�f���;>�'��؇>�FZ%õ��L;MU���ψ3�lG:�fe�NP`�tB2u%����'�I����&$��11_��������2$��u�*XQ�½�����fR7);ܫJ�C��{]Zl���h�u�1�����-������I�k���E�u��ZxX|^N����t��Ɵ��^���$���"&%�Y�o�b����wU3g���jA|�r� ���E�v��=���i�>U���^�c|.f"U2�h��5��ҏ�T�l��C}u	�[����/�;B��;H:�^����`�t�%����^�;��{}w݅z��b��d]{����ע�9( `i>#�ϕ|/|=��KJ0�?x���df,�B¹�ztx}�C��7�����Y�;���|M�k�925�;���<h�wxBz�	$��!�&J���l�
(�R��NwO���O
�k����u��<,>:I�{~��b�����4e���+��ʻ)�.��)s\�f�*j��гCW�����ҕʔJ%H��E�J:���i��Ua�E�֪�a���s���]5b���<�K�ũ6�V�'Sӣâ>����N� V2^4Xm�}5��̮��Q���V�-9$2�/X�7�YyP�Çr^$�<`�?g�V,(��ګE�fN�vsO3��i������bw��<�91�9�t�02�뻊�A����)i-�o���
n���cz��|/�|�jE}w A@a$BaW�@�ҢnS�<��>��	���C���rD�1O!c�h���|��񻬈:U��'�n���B�{�}�����τ�&u���T�*���m��w���q-B�W�_Y� ��[����A���m$Yi��I0��x���w▞0����h�s֔h�3��=i�a�vw��Q̛��#�JJ�F�-�ô�ј1�Z�+�������p�s)�g�=��94���t(v���Rf^��4�Y���������E�7�$)-�x��KH4�|��<:�u1.D�a��9��Zs!�H�!�9fl��h�iC�n���
�>�ĲI�zD�OC�O�K۝�UV������x���~����2C`�-,^����M�g��aB�é�s_\n8a����ty���  r}�e/�4�ܫ	0T>�V�,92#����PϾ�Y�g�ؕ�LJ���x��ZA��ʝ��L�ܚ��3{~ފ�E����8(,���b�g�"��*���*� �
 ��
 ���(� �
�� U��(����
��C��%`HYBF�� `IBP��!`Ie�%XBP��$eP� HP��%%	HFP�`HB��!�%	B � 	B��!P��%	B�%	H��!�! HYB�%	@�%�% IYB�� `I�%B��%`HYBD�%%H@�%`IIBXRP��!`IBP� H	B@�%%	P��$IBV�� FP� IBV��!%X@�$`IYB� eHRP��$	BV��  IRP��$e	P��$e��%RP��$%XP��  � P� H	B@�%%	��$`HIB��!`IB��! IBV��!�%�% IB�P��!% �  HHP� H	BV��%P�� eXP��$%	H��%`HYBB�� `H	B��%�$%	��$ IBB��%%	YBB��!�%�!FP�� eHFP��%P�� %	�$%HRP�� %��! HIB��  I`IIB��! HBB��$ HB��% HIB��%eHP��%%BP��!%	XP�� e��!�$P��$�  HBB��% I	B��!� %B��$e	P��%%	H�% H%	HRP�� e@�  IH� `H%	IB��! H	B��  HB�P��!�! HIBR�P���! I%YB@�!eHR�%	IBB��$`H	B��$BP��%B�%	`IIBB��%�!eBP��%%	HIBB��$�"��%�!�!�%� `HYB�P�� %	�%�$ I�!�  I%	BR�� `H	BR�P��%%P���%%	P�� %	�P��!%HP���%�%�$�!�$%	`I	BHYB��% HYB��$ I%	`HH	BB�BYB��!�!eBP��P��  I%	`HIBHB�BB�P� IIBB�P�� `IIBB��  IIBBB��%�$�! H%	BHRP��!�$BP��P��$%X	BP��� %`H	B��&�P���&�P��$�  I`I% I%	P��	 HBYBYB�P��!� �%�"P��P��P���$ H%`HIBBB�P���$�!%HYBHP���!�%�!%	� � `Ie`H%	H%`H	BP��&�� �%%	`H� �%�&��%�!�&�P�� �$�$ I%	P��$�&�P��$�&��  He	`HYBP��BA���!�$FP��$%H@�$eB�P�� 	B�$%B�%	�%XP� IYBF� HB�!	B� IB�$IB� %B��!P�`H�%P�!P� I	B�!e�%	�$� `HXA�!FP�`HBP���% HYBF��!@� `HB��%`HBP� IYBV��! HYB�!	B�%	P�`H�� @�$`IP�� B� e	��$P� I��!�%P��!%	XRP��$	B�!e	H �!H�%X�%`HP��%	�%X�!D�%`HXP�%`HBP�� IBB�%��!`IP� IP� HB�$`HP��$	BB��! IBP� IB�$e	� F��% HYB�%	P� `IP��%%	��% IYBD� `I	B��! HP��$e	XP��$	BD�$%B� HYBR�%HP�� 	BF��!`I	BHFP� IBB��!	B �!	BR��!H�P^ �
�� U�
 ��(��W� �
�� U��(��A@�
 �� �
� �
��b��L��51�+� � ����~W�@���į00   t  �  @�z � :  �h     @  ��     .�                
          P �      
�                                  @      2 {��R�=�A��79�4���S[��x���� �v�C=�q*������-.Yv�P��t�����z��ًy�톊k��:T(   |��ϷG�4�^{Pꔛ�s�n��ztz+���N[f��z�/0 t��� �;��y�^&�{����8�u��lۗ
� F�      >@ g{lѓM�ƺ�@�F���.��F^���sYK� CNؠ������G�� �lQsztW����]n �{��;c�a�h�9�Z+@@��C���:(�;;f�٣ g)��+�;�k#��n�OLA��u�ݍj]�w��mi�-�� wt�M1�Ľ��v/,WZ�7]4Z8��҂ �  �  @    ��c���V�׮�=�8�Qsu�E1h�΀������i��#Kf����B1����6́� �i��*ng{aأ�hu  ��(����-=�w��Z�C�إr��J{cy�P���3��Q����zogC7���z� v�.\W���[�t���=إ��� ( �  @  �.]�٢�������9��f�4��뢊+�[� ���9خ'�:<��i�Mv�4�7.��  t^��owy��`@ 4w�נzi����(r� ;=A��tz/1����(A����p ;���)r�yV�lqb�E����qٻ�y��C�   �  �      :�ހy�w�tQO䋠sn��C��r�R��&��st�r�K�C���p �]�Nn�b 70�  
H���5��y� z�� sC�=!�zP��׋�y���6{��֍�� M�E�l�=H��x#��AO�   S���J�   h  "���4��P       � �!M4��M���z���z#i��j��P
UP  ����� �?iU=OP 4     i�R�D�=@h    �>�[�@���/a�ӷ[�7κ�k���|i��q{���UTm�k�EAW��A��*���j������[��~X??_��눇�PU�Um�b�����0�G�δ�5�Bt�m_o���?}�\����i��;nű��b�K�H� j�� J'W&\J�S�C����VVu3��X;�3t\�S��nf�x�VmFS�{�Qî4+Gfu��)fw�lɈi�"�:N[y��]�n���q��7�%��U�bU",��\ݬ̫gC�
wXw���@`(����w���l��J-�7V�V�wG0n�u�i�[�����6KO �64��w%�ױ�q��3��A���[������&���ѻ�5�A`7D 1��ɵ??ȶ��;{�kQ�N,Gt=�sv��̧}�b�\:霬Df5�s�e��O�ݩQ-"�,eyB��wE�Q�(�ͣNjf]&k����Z�����R��p-̛oF㈝ɣ6�diUᵺ�n�a2��X�6��>����Mf]��GX�偷h��r=*�ݱ/,���]qO��6���ନ%�̸��;:����Q;I63c�,�Uxcy#�sQן��y7j�piVI!���-�����k\ա���V�~�t7�P8h�n@A��QlW@6��hZ0i,�Т�m���F�]�B��l�ݷlm��}��Vea��)���y��˥��Ie]�kXv��1�,��n�Ƚ�%����X���������w~�\r�櫹��lu���(M@RэaK�"��3�ٷ7&���0]�4�wj
�Z�Q�'��-�8����J-������\0m��B�R�;�ŉI��ql����N�-�^̚�b���������j����� ��qJ/^��ͺʻVy��~n\W�f��sp��VnΰjJ��p=�u�:c�(��w`�ͧO2�N�b8�[WfTE�@�I��۠�
GE�Ɏ7��J���RXgS�!X��ZCC�t2d�Os4mn!x���m[0h8�����i~ܲ��E*�R�/�J-�9��#�wY����@x6�M��o��а��ʭ��RBRd��Ak���	��S:*�+R� ���U�Z�e��B�¯oo�(��l�V	�p~x��7�Fa.	���*�N����Pچ���t&���.��v� KV[��B�K�B�Uk�ܼ76���@D�NV]����q6�� �p�-鴶��T.�.�R�PC�U]�ΌP�	�Bn<54m]��^ӎ�4�f�w�]j�ˇh曹�T;/E�0U����ql�5����E�iGU1cՀ����jUX���ᚲ7z��x�*��2�i�&;��U�M�V�Z�m"�Yf�2�`�9�(���=�X�Iڦ�����$�Fw��ь��c����ț٤�֒6`&�[��� �&��;4ӂ�f�ڛ�f�BjWSu�7Wuc@;X��FbpeL	�7p��e=7yB���͎����Y��-o5A���U���%j4�ͬY�2�`6�zq��ݨ詎��4e�l���s@��]�S�j�hp��N�fV��.��&��VVe8l�5gEjcq���g��u���w�ǖ�$���ZY�@���.�!��,��Cq
B��[�jZ�@�f�2�Z��v�w���l�ܓ-e��mm���VKr��LV�ǧ/Ue�oul����P�ND�,��{A�ͷ�cT������RSi]4�{�h�/j�R,hgS����8k�&fӠ�`Շ]��
ѓo*�5�ʕ�#�<��M�Ij<�`N�雙��6��"�d�A�4!M���;ln"�g:�fT������d)Em7u2ݕ�L��QX�-�U���L�t�:?7��ȵV��4�i�M�k�J���үd�6�Ƶ,�CYFe���{�ݝ�R�׆Rs�*�,N#��g�"oym�=�	�B[sj���a�F�y�/"���t�{ub��E���]1
�/j�TYW�����;B�:�-�x�gb���F�;*cJЭ{�ZE�yY���m�?�5Xl�SJ/�3I�cw/+m]]�N�(��k�kR�*{۵J��iJ"G��y��4f���C	��i�l�nk��T�Z�e�LL��T$�i۽�w8��b	�a��<��ooX�L��v�y@[5w��z�ͧ6Y�B�m��.�_e���!X���< ����*h���ܕ{VH1��n�j*��߮�U;.�������n���A%n���u7e�bg��3,(t�XWucp�W�wwd�[Ki����֛�
�X�
cf,���Ӈ4����,��(�osHC"���w�*�d0^�֔�`��G?C�tVRFU�c�u%qګx"���\ۥ�LX��B��kwipK��6%�M�CM�LWwV�cvm��fV&*XETLf�XǶ�P���.��uP��u��tյlO*Ŕٷxaʽ.87s*+;-��8R��L�V	D��f=���M2�/[��[Z�oavImց��kٚ����oq
yQ�pT���S\�8(3	��D�+Y������4沔N�\�#�U�ri��f6���#W�@�ͣ{��F,����vnS5hīS~P�܃w.@��������f��&۱z��$3+%�����C
V����)���;�:�m<�yK-�`%�oH&+ǦԳ��Kv, ��me
kh�!��bx�!�%AR���P���ŏ3u�FV��b����Vjm�o̫��{��K�`T�(=����,Ѵ�3TS��oL��R8�o/!f���9{�4�J$L�R����1�ݼ�B{y��7�f����m2�'��Hp`�-�-�<&�T@�ff;f�hU���!U�/C����D԰o:����e�i�2�������4H�e�ݰr���R��bv��ʔ�-cӷD�e�����m�%cku)$���-�٬�ʻ��]<��f#7B3hF7]��J*+3sr��2�SZZ�e��cvIE�V�^��(��jZݱ/D�{��*M��r(g�6�d��V֧jݲU�M�c�����4�V�����k/]ГP����s2��5�Y[I�i����s����i�^Jۂ�i�5�k "���;�z�e0��@�:n�Q�,��f�|���= g��YO/)Ҿ�8s��
y,ѣi0U��ۙ�W�.<�M��b�Ck5��x�օ���X�0k/elqڰ��V �k�Gg�8k#��[z��a�w73�2�{Cim(6T�[lӐ�aXt�j��wY5E�c{�D	���x�q��ɢ��FK�1�U1����.�15l�id�Wkր����X0��O-�8 ���R��5��nf�����&Y*\�����V���)��F��WOK���V^��`�۹{�r�fP���nb��d85]��0�3�0��=N�֗W��Sn%�cˬ�/ {�(V��K����6��'F�ؕ�T��l��[&Vb,��Ue��Z� �@x�ߺ��!�nP�g�-��I��.��V�!�H֙��64QըT?��y�x�ӡ--�2�a���-�N�_��]�Jj�G���W26��)B�em˭�T��������BƉ7A�v*����] m�CF����)�z�� ,K#;b�û�]#�
�$J�/r���b8S'//6V��RK�%�PSSѳӟ���0B��l��B���k2m
נl�A!�x���%䭻����/*Ł�j6��,e]�8IO��_�#Ic5��ZM�տ��v F��(��"V�Z��[t��N��)n���%n'NbJei���ۢ���)L8�ƈ�i�*������yVͺZMӖ�ІZ�5�S�I�P����� d/k�Y��٫U���1?����A�1���p��Z��7�6�+m�9*f�+ <���^�2��[{��j�^�N�1P0T�KvcU��[�ݒ��K&˺�i��R��OeDbx^G��3fc��h�i���$��P�ב,�ݹ(��k[�կiH�3v��.�47����Kiа������or�j��(��p��
e�`�jQ7S1iI{u�XYsv�Up��Q×Q�7�t*�A.�ȸ��#��b7�	�8<ęp�f�VQǺeG�Q£�T�-^
�X�]]m/#��e���i��b�%��y�Pw7nM��J�7�J�?��eC�8[���l;Q��`��z�V��cT�`�{GE5gh�6%�564�xKq��0s�u6���"��Q��Y.�2
K.c�(�sA$��rICK�{$���ST�y�F�LPِ�rΐ2+3@��3n��m�eܣzn�8&�'�B��a�� h�$�/n��B`e��.����R�H��Sʇb��I(��+C+%O0f��n��6V�w��-���Z���Ve1���P�H
�����J�[�e�UN�3�:��I�n^�Z�fB�tASN�i�BEqM!X`� ��(�S/%���2�7�`ѧt&	ܽ�eY�i���L��kf��kg�d�<�D�j�7.��jȚmO�N�F~9L32�	Ha�wXwpǙ���a`"�fE[�qTmQ� � �+^�ٸ��j�ޞ�P�������A?������T�4��ýn����t��[��+	bݖ�f�qݵj�����҇C�j�LE*�ܛY���Z�e�]�%nݼgb��Y���b{�5�,	��$�kA��2ɩOu����#S5�v���fQ��������`��.C%,�2싽����M՜��4�V�嫙���6`���9�ׯMn#�i�1�.m+lu���^����w*�f[���[+f�k������SF�{�-R��	��MfT�˹�&�m��ܲFMR(��S6Y�ss/6�j'��z�����R��cY@��u�7&�<&ŷR���ee$^V� �WR���f�r�"��鰣���X����L��F��j=V�L��R��F��[.�e0/7�o2���e]�fK��ǚ��Zr��c)�+��먮��Wᙙ|��{f��ԍo`�1MI������dMǙo,�bTD풷?]���ݭ�gE��nE[������5Asq�M�ke�ZT��7��
���޻&Νg2�ƴ��m9��˲nn��\�7m��Y�x-��#b�5���p��X&��c�yI������,L8K����f=�w{R��c&�͙q<�g��b��RF�F!&]��G(ǩ{VJn8�+�n��E�W��ѓ��lu6�F�c4uیmּ�Y�W��Ǒw,!Y�T�EX�vB7�QF����^d���k׷���Cy��;r��e��FX��aU�е4��f:�Tj�^nb�jeC�Y B�n�c*��]ᐭ�v��#��N��y/�s3q�{E*���n�J�h7t1�i�F�M�:��!׈����Y��d$��rj�����q�;�u�M�-eIBVh�N�Q�X�:eQq�Ԏ�b�Ӄ,$D�y�&7ɚ��V�o] ?H�*�$,M���АZ!�G#ʳqRkZ����l��d�;�3*�7&f֑�_^ݐ*����"&��<&�*����h��	�a�UekD����G�gB��f���!ˎ܃�Y�)�x�"^J�Yh���4]�:n���$��t��$1mc�/��ޕ�W[�t�&)����^\�ZX�w�����[�C2�.��^ܑf���K��c#�U{4�_�u,�����b��6~cE"�i�G/
Ò�=Ĕx���@��mY��A;�{���AA��+(���1OwK7z�(�lba#7t�HJAV_�[�S��䡽ֱd���
���f�c.�s
�%J{�Ѣ��4m�GᕶE��2�=���{�B�V�lȓ�Z)�I��������(d�iH����xQ�2V�r���C34�����Ǆ�9�l�����R��v�W)�T���^ݹ�+{pZ�0��zB�lأ�z����6G�xrb���y��� ~iچ���c-q��U�fG�Z	k^�������*��X%����Ts��e'�l����zQu�^F�33
[�-�u]n����5GJB��[[�+��%:��%�TNE�\Y��ZNcȳv95��5��TP)ED�"6sM��k)��f�^%�Jx�������R �4jKg<ZE�4�V��Tg����MV��V�O!��n#�n�V�&f���r��".��8R�Mݱ����[4�4��Ɲ��?'aM ��6~v��������T���%f�{��#`s,O�b�[��m��8����X��ԛ�fE��U`�.��rKۺim�D��fSnB6�VC��c��2R7��y{�ջ��mQ:����J)R��� �0�k-�J�@ʻsVmFu�3z7i����U*͏(�AK̲e��&I*Ɩ˖��.�97niP`�(̈́�`� �OC�����܅���y�3�47�" ����&��;f)V�H3��� ���Z3��b�*�.�e��u���n���
�n��1U4Bu�ܗ�SBe,��Ë,�mdkHЦV�Py�'yd��+r�9qK�y�	��x����nnV꣔���u^���E��bM��[�ӧ�S��ՉV��X9S�u�C��]�����m��Kaf�iOH�­T���0����۫�M6+6o�{��-��Ժ����P-"�ғk*�cN<Iy�R�-�ݭ-�ق� �KfI��Jǅ�Rn=mv�0h�y�3]ۣ�u�`:�(�3/e<5��.�z��bUѦn�u{��`Q�7^n-��� �G]k�n��4X���c�GE���3c-��e��3BG�r�3r٤&�SUD�l�-C+���ckVo���hG�@ZHxhŹC-�)n�)[�U��xsU]d˂�I�m�!��Uب��j#n�T��4�ѕ�e��,�ʣWl�����ԖXa���eV�F�rYy��(l�q�5�ܥ\y?�c����T	iS�1n]"l�*ȵ�x��kcv�[xTmL�}z�e�L��'wI}�@�@�/*Lv��Ю�e�� ź½Ս�ej��a��Vw_*���ۋ)�{旎���6p2��#{��ͤ�3��+�Q��J9�u
��mw]IrcwT���f�Xb�1�]?~>�_�~���ߟ,���
0 m����X:Ҥ��X� �[+j�-���[������rb�Mqv�Ấ�ʬf҈cl\��cip�U�������̺X�0�ٌ�Jj62��j��X�	��(k���)4���%���iA+��������i��j/	e����X�X	���\�f��.���ٲ�ؠ/�C�ᕩ/��]��t�AK%6�
��[
I�_k'��Xum�����k�źGVKdkMt�M�`̫s678#��rk�])�26X�'v��J�ز(Y�4)ԙi)��ٱ�q�l��2��1��v�m�m�.�ij�m��і�3IJ��[+�ս5�Q50ic�f8�R����H����Z�&�m�m�Ąd��7Ky�i�ە�^��\]2bhܶї��gU҆mԴ��n�hQІ츌銳XR�=V8ai-�5��F�lj������U��(�,���:X���u��e��u�+�e]��q	���e������x<]t�5Ýw1C��i؍!�!�)Cj:��ei,1�`EMV��ͩ�f�c���h�qm��36�`�L١�\՗L+��Ku��R޶$��]��ԉ�ˍ
�7b�ZCif!�X�Gj���F���c��e�kmKq��ْ�e�M����r, h[ID�k����Wb����[eYc����[5ԡ�CV�R�h�m��0[�K�i�u�6�J��.��]��^�HL+u�7hو��i�K��
�3L����4Pu��6�[��It��pM6(m+;f6�͐�m�\:6X;-!G��]).$���4%y5u��۵������T��j�֪���3��Mcq��k�)����ir�9%/jk-��#K.4;n�Cic�f�b���B�l�m��B�l�喗i�P3ec����.���]]�܅��[u��k0J&K��sn�һ���f)LK��Ʈ���
�Q9�('iY$E�2��h7�e��kcه%�ZK.�Y�sm�������Ց��M��6l��Mz�1JF�lˣ��E��Sҧ6Yu4V��*�m&v����fi�cb�v��f��s
ZGE(���ZbK����W�]�]tj��4�n��J�l�+2�ō ���Y�b^СZ�u�%l.̔��[K�kL���EwZ�e�׶�;�IH�	m�`����v���ۃPm�t���c�n�i��Y�۵��.�auKK��cqc�l���ؚ 5xK�WRl�ڸ��b�066�U��I\��j�klM��E������s�帶����X3]�b��I�����^�m�.fs&j-�j]Xښ��V^�az�sm�$-��S7F��R�E�\vi+B�1����� �MGkV�6�����z�R]-ئQ�h�����X$RX%ԭ[))�E�[�jM���v�X�S[Yn/���mɃ^�Bl\3GZjL^FmQɬRe���|{�8��]���H�6P5�s��nJ:�2Л�׳���I�nE�]pm*�MIl�^�q������]:�t#Xvc]��K(k�2�ؽ���6������%�j�[ݬ]��\��U3Z��f��`���s��V���+Xe�\#v���}��Z����h^&���]e����0Wq/mWbh�YhT��фm�m�$�M/�.h�)ly�����B5n��u��6����@�m�S��TdH�ٓmv���"��pèۣ�F<դa�n�b�:f���-�e�6���N��*�P@�3KV�Q�F�A4а{[�$�M��K�#�g#�5n�i�J���av��X���CM�T��ζ�t�YiYq,���H�V���}����KKn[lv�,V�Hl��Z̵���u�ҥ��-(�1��v���iH묹�6SMu�u���n�rJ��MV��Z��֍ai�S�$m��k����6J�M6K�b^���em4�t�XR�+A�5��1�4e&$5��P����m���.����@�m.��L��t��������<�[p2�@�m�G$�mju���×_���_6mn�T6&�;RIxź6Eًmץ�eeG[!�ݠSK֖Ycsa6]��w+1Ji�
M���)�٦�Qp�Ԁ�e����6��tf�P��8�5���C.VĆ�B�v�M-<K��bU�Zbn�m�\���!���Ͷ��ҷU�j��kf�sqԸ�xM�����3MȷF��і)���e��8�jc�bP�#���ɋkM�:٭Ѧ��P�Δ����i-ʐ����5��q�la�JmrYIh��m�mI�����V`ל�k�1�;h.�8�
b��naJWjL�č�kR��M��Qq�����.�,��g[E���eΰ4�ˀ����\Uv{b2�[s�X�*5x�n�X�K�=h2�Mv~o`��k�6u��Z�G�ͣЪ�`�Z��vL�j�Wm��	�B4R���*�h�R�Ҏ-�L�])-��҆�0�mMC�k��[a�d��C+��iX]���i���!��H۫+�ڃ�\Fз�#`�H@�T����R���-N�b�4aP!Rb�K�h�v�9&v�L�6�V�P�����a��6�mf��f+��:ŌΤ�壍�ƀ�4K�Ҍ�&{�ۑ����ҹXk,�:�wWz��b�65�Q�R�M45c)��M�8��d���	n��ZZ�m���iN���I�,e�4�f��-���bʹG��./�=c���][]U[�E֡�
��0��[�ʹ��Si���Mk���؛X;]��M6�6�f:�VU-j��4����6̤x�j	t��ˮ�������e*��у@��cJG��k�-,��#�lj�,��Z�	j��-��9�k��b�f��.Ê��\�3Xk�v�KoR���i�#e���([leŤ�Bݫ�+v��d6��nڨ�l�2�ؖj��NJ���m�a`���a���V��z�+�vJ����!�F���\֏^�v������&,��&!-���CB㫲�e&�%٘��5B$���]�\U٢��V̩3f��6Ǝn��pkm�K�#�4���-�"lӥv��%c��,ױ� ����v�r�l�kb5��i����rY,���AXf����5�[�Է���0�n .қ4�f]av�ڔv�C[��]�Aٺ�[BKpBEc�śM�X���D��� F]�&l�M��k�KMs,��KS#�MCv
k��jQulծ��F4���Ne���!3��J�)	tS.�qatg����v�B4����m.�͊�{������Bvڮ�3l��lPs���e.�K�s<�}�fت��]n���T%y6[0F��i���u�a� �8I��a�&����2R��c=m&��%qZ��`k*b�n�-�ԴN-!e�8bM�sm�y�q��
;�ʵ�z�&�%oX�)�k�P֥�e�S�k,�Ѻ���1�bM�k�s�m�nh-��-+͇j�a&�l������[�ʄsnŶ���4�-�Zʷ#�4��%����9��L�;biH�X]^��i��9�����f�a�����ԀKCp��F0ɬäil[fKcV�F�6�`Qƴ�0]�3.��DB��0�3�q.[�,v�(L�kt!��b�ZpTM(�#v;iZ
m�]�hnd.�.��]%�@���i�y1���,��씍��J͵�7b�[r!KTv�ݥ��b�U��M��i@�63v��C����8��!4�s�j�ݳ-	E&��\;���x�]L�fՌrF2ƭ�tV�c�=q�8��ж�n����l��m���4��.����[X�Ѻm	�Xd��]�Is�Ђ�oe�[4��,ή�-k1�u#V�g�hk�&�����vst+���b��Yup�ΔB�z�*ٯdl�(MA3�a�j�����b���ۭv�.��D�R˪����k(��Uj�	� ��0�b��Cm��jja+Ŕ�]{,�b[�[��L�L�p��e�j�0]����A���k�BJ��m-&�`�P�f�K6��pM-�f�4K�YV�B�n�Z�GKM��j�Quuɶ��q��jꙍ�RQ�\��F"94MB�Dr�%]`�R��h@6m�������&�2��_�x�M�_�)�g����M��+�n�TAƻ@�iI��kK5�����~`��:KGF�|+,�SW@�Y��>���P֝�,45�e`KRW�:�r���XL�QiM�Z������i�n٬����h�-�f��]@�4[nv���һk(���4,4H�B��,�(6 ^#��n� Lk6�����\�-Xnq.c5���͉��R�M�v�FjF0�Һ�b���t�Ѵ�m�Ɉ��5�j˝Csn��e�f
Gk�8&3j��̻<l��������Y��V��1��M���ٗ���\���:Z�2����lݙ�Rl�:�K�.���Crl��j&і̹����S:fb�rR労,bmk1F��F
D���j��l�gLm��1cl��ܚk�5�F���<)�39�W�i
�iu*\�Ħ�qf,�m��:�R����s"��$n���͛��mR���L�a�$��,aJ���f�B�mɢRR��؅��WHGiff�f�06�mQ�z�1�Ҧ՗D靡KJ�v�J��;�v-dt��e�%�F�s�N�醶L��.�^��-�νn*��b1f�٪7-��̺���S/P�&MY�m�L0��E��Bۧ׷^d�o�{��l��kvY[6$�x��&�+�`͈��om4�m`f�n��6/g�2[��.c��`saqpM�@u ��rǌ����H��`&u����4*v�
�l�����T��ۣF�QqV3Ԏ
�&�f�:�j�U8�].��#6]f�c]��\:�Y����2Q]Kkh�3M,^��a	�d�< C<)y�%����=j2�f�"���c�=�H��JO]vbA��M����摤ɴf����R�	aT�Ca�a-QZ�����kvt����^����
̦�8��a��h����^&ųE�Tc�a.2鍣HY��[cv���0;p�[sa��F�m7Vf��timkK�3ےe.�.��g7�k����etك-����h⚚��@��б�n²�~-��v�9�+Z:Z�!&.�)�l�K�F�fM�V�v�s��Sh[Wj7gB�%�t9L�%c�ZX��i�Kh���mn���4�M4t�&���541Lk��X��5��%�6�@��ha�Z����U� *���� ��契��3�r�թT�F�ѩ ZD� B~��b�9�YW�Z� R�Bc�E�K!��@�p� Q�:��Da����X�pB !�# "� L��:0���/�@8��,H�x����`C�$��	&;T:,x9"D`pB�@��*� �����H�Ñ# �2�B4���@�b[�1�?�ހ6�(T!*�*��+�hD�e�a�DP�m�E�B�Ycl��
�*G�l� �@���c��e/b�p�p�V�D�m�%*�"�!�#(k�+#�bȜŏ�>��^ G�@`đ���@2�$��f��Z�m�!�僁*'��Ad!p[Ie���/3IKal�N
,�a���ґ����C��D�Ͱ�b/�-�E�#(�acFF+��Vx^X�� p1D�8��,���+ʤm��X1e-0�ң3ԗ4�V$5B\�
��GR����$D8�Q8�
JX[j�^a��5�R��$a�����	/V[��` �Nnd� �NC�[/IV`J�V�,:�!��)IKh�0 �f�{	J#%�y�2�X��8��F�b"+2�!ʑA!0A$X�qil�LLS�V�1�kJ�� @b�" =������9�ƌN �<�p�>�X���\�Dbr��:��
�������T�UN�R6�U���$8�\M �� ��+ ��o5�U��Jup�ס�,9+��f����- �n�k�%�bl�H��N!�U�[%�B�
�m�HA(�
r��H1!�j�J@���ZS��(,x��G��T8y9^EHD�3��g���/"a��O���)X
�kN�J�Z��-�R�II�Y���^D\�@Y�S�b��*p8J�z1bmf��Z��/AAP��。�),�k��x��F*� 
H1� @�����#�	��(�q-�Y�,I�@V	%,"R�NN��H�B9!bJޱb@z�	�P�8��*�H�"ǡX�րrD���8��@����V�0IQ� (� G���Kʉ�n��RrI�JK ���m��P�Ae8m�-�^�mT� o�YMZ!*�@���
��� ��/5B!�?bB�İ�*�C��(�Z$�&c 8�Dż�������"$U����@DYJ�-��, #!BHE<��' �^	(VX�1!+V�Iy X��y:,��m��)���)z1m�!DKʅ�����K! v Ls�� ��!�,X{��8��"�rE�1B�����ǧ�⚱�e �c�B�ÒR�[l��KP��$AF1N�5�E %:�'R�E$+��B(�XV�
�`*H�dHV`�a$ NNH�����H��8*�RZ@�pJs�#�$B G�c[^�/t[JimJ�"� �),�x�H��o�J�R���C��$t*����Èa-�x��%��E/X�y!��e���DC6��D5�Ŝ���N�3�B�@U%�Vz����J��H��^�d�q��A�,$��,V�+%# HHԲ����$p$V�Iyz2�5�Z#��A������c� ��a�INaQ�%�� �y8V+�egXS�d�= b���Io0��<����	���R��^8��1�#����� [u8����@1iqã)�!e��%�-�Na' DQD���D8T�@"�4�S������e^B5�A���1�z�Ia+�#�Xŭ�m�y����c��Ԅ���H�Yi[Y"��;�' t�XW�O��! ��!�pr!��	�ud�5 �8�I���J#�e,) �Č*6���V���^YjI��XB���JIk"[e��%�D @� Ùȁ#�d!���C����2�!V ����0� �q�D�NPa��\�
�e)`U�a!+-S�H�`!akKP�K�� �R#*�D&e>���Y�HIH��!B�Hp�q �C� W�U��# T	�)D�;$h��"	"1-/K�KR�J,�e�����}}�9@��1�X1� EiD�9��H�D@x��-���t 0VD�	Ā��Å���"+ehEA^e׶ ���I�F��B��'6��5��XB ��x!:f!�!� � �H�F ����b��!:���V(p��[z� �o1�!�S��$$�y:�0a�E�ND��#+�S�1$�Z���B pTx�F,U"0� @ Da�8�^N%�1�pC�<tel�G�� �"kR0D+,� rJH��',c��bD�q#kcE@X�/pS��G�ǁ�}P�H�1N@��'D ���J%P�F�����P����R�PBXx�*��=b$"'B"p�� Q� �iA�H�	^':�!`��F����(Dd9:,^�i(P�&�!"���bp��j� @����m:4�D�J�C�V	Ad"Ø��� S�ŗ�P�2��R����E!*1X��!��N�Bd`�A#ē0#F)6�z��Hpr�֐"1c��q @N$I2Ł*��� �����6�iB!����8��G�E�5�X+� $dI~,�����jB6*��-X�� ��)T�BC�Ȉ5��!� D��@�3�Ma�!�:����<N�[V������8�  �(�F9YKP��$ �X����89Ug��n���B+ 0H xHBu���I��c���&�y@-����,&y�!���䄭[FY	��
��I Db��Y��*"A$W�C�ef�BR@IC�����"'�g�kaE�r"D�@ 
�� �<	 �x�а�"��)<�rD��b�� yH���/=H��O� �HB/sX
�Ъw )ޭ�I�� ��$�Y^H,`rFQ�x	�FB9�^��ʜ��p��X��1 )H�<��v#�I���ǉ(ã�R0�v��� �'sdFV`[�XB@��$@���P�@# 1��p��?2x�� ��K"Q��JP9�E�pwé/p�$88�y*�H�6�q	(�D��EW��8��Pz�QN ド	�	�N F*HÊ[�� Hp�UEb�����<�F�B��(� 
ʧPeiהT��
�/"01��z� B�"�:	T�d$��%�d8㭽R �OF�"tH@^`z�����E� aH��!$g���Y��n%1kH�!!�a�w!dB(� E�)s@�W���<'$�I�C�bq +��Ã�a�G��ˣʴ�����F@!�V*wAx[Y
ǀ�H���cI�H��db����8!	!	"ǖ0�3�("�q 8� �	 q8�R$ �"0�"�X�P��x# �2�YB	>Vv۴R�!!:��@���E�
�bJ�X�k%��J�ԑ$NW�!F�QXJp�XÎaҶ��  �TA�K̈HD�@ u#D�C4���J�t��%-�		B� �#$!�,����Lǩ�)��	  +��*
,��!	D%��PZҰ$ �PG�u)`AH�Q���YW��$D���B!<�$H���!�P��"�"0�X�@�`0` @�q+̄� �N��A�,�$c�#��<ʨ�J$��X=���� "��Ėtډ�! ##�j�R����"��jP�^`8� �B,�)b0N�u���ăP(�R0���z's �F���qx& J �	��PA�� ��sԫ�1$�+� �3�����^ �F�S�Ai�߅��a>��0�+�$H���1��(���,R< Eb�`�!� @ġeR� �V �bH�H�!
�A "0�<q��H��KUC�:� G��*� W��d�p0�ã�H��ED�@/��tN�!^�H4�� "r#B�PHB1���ey K8�KP�Ľ	۞0�J[�t �yJ�Bb�a :�"�B�b*H���%�X	���Z�$�J�$ ��RFR0��V�u��P<���-l�
�;�=�&� �(��� �@�<r'r1"U��$!�BEgIt �D�  $�EX$�(��O�q�$E�m���ՈB  $JR��"HC�H6�t�!!wV�NH�b! �@�$x��# �Q�<"H�@���Ea��?���ù;��r�P:8"Bc  ��Q�0���'$D ��'�X��1C���I$��AY�l�@�im�Z���{�(�jN��T�8�P\#h;��%]���0�+��*������v�����0��f��-6��f��-��V�bX�F��5�M+5U�܊�i�P5y�V2����Ҷ��ˌ�LֳY���&͸v�!��.Mu�69������+&[�6��s�E�#t`�\�����Y�f��tk���v�eK���j֢��ee�lqn��4q\gZ`���b�Mű�SR�6���\���i56wP���[v��U%GF�be����#��qf,e�ѳJ��+kZ]j&��ꁍ�RVlCm4-iv�b��u��Y��v����Z�j�x��;k����:�#E	�,�Ɇ&�n.P��m	Mq��RSv���]4�ٖʁM5�(M��	��bCAJ�CHm tҰ��jL�ِ��m23KR^W�l[�p��m�V	�LB�d�i�[[j�!�r�bgK]ZJ�&��jE�M,5�	��.��{m�B�Cgbiqf���`X�Bn��=����rۭ1�w�%c�V�M�%�R:]pǫe]��œ!4f+ L���!mv�Z���a�'0���\U�s���rį������p�,А�Iu0;j�F�!0)��5)-��i��Ks-�L:��5�BҬ�bY�3��d�L @Xa!(R�${Li��XdҲ��insm�)�,m#G[W���e�Z7i�MeRf��i�t\ljs���X^5��c	Fͭ���&�ɱCiP�m.���݋��M0Kt���-bK�fq��2ke�l�v�
��m�m�C.������QKZ�͐�K.��jS�m*�%��+���f�mڬu�.��0��M��e�L�D�W]4L�Sb�Ir���b�Kvm홒iF�ܙ�j6��ѷ.���P����X[��v�n!E�\�]�M�غ���M����D6�@魃�]��\۫K�\��JRB�����Ѽm���S� ��UKe[���j5J��Ѷ` )-"w���)~d�T�1B���Q�+-�K��l\�Ui��s��m��:d�X�k�M�5nn)��@�P�F�
�����x��Z
#d]3|��6mݮ �f]f�6��A�1vLT�9�j���КZf%�cZ]m�a��� ��V�Zmn̹���Cd	�Pa4K0Ú؃ZF��y����fk�In��F�E�n�j��cb��-�5s���i���ڀD+����3uUŁ�����wl��jKi ڙ(8��e�[e.�N)�<]^,�m%��P���e��;P^��.��Y����%��-�H�#mloD--�Rƈ�šR�6TK�C�iT��Pm��wV�[���i���g2^��eM�J�#�o*����g�=q�`����f�93�����4]���p�U���^�W�������V��B�+a���-���&$�S�	�)�=u��Λc�!�;�����r���'�=�q�\�����ܐ�R�'+h�*Iʹ1;��5Tu½�����}5m
v����a�ֳ�sVen٘�!O.��5�����F�?�@*���V��� ~tM��@�9����fdV��j
ʏic��O;6�6W�;�0ݶf��U�D�i��a(H�a�i�H��[0*��|���Vg�)ŉO*ujVw.M��~8�_w�s��Աk���s^�0�s�D踷��2���j����W``�8�K-ݛ�m�gB1���m�ufe�ia�QJ;}J�V���@���2���º�̞��P���ތQ>�9��v�S�s~�T�������]/[����y�2� i�Ji�}1t�{�z+7� q��z�>���۝]��l�UL���V1n��5���A�,j@R���5T6�v�ӛ����-�zX�\���ƪ]�9��������:��;z1n��'��w|��I�T�6��޻վ*�g�;ݷ)E[�1R83��͟V�:�btn���7^�p���� ]�M{<)��"Y�6�\��˙ݚ�z���9��nEed�(w��3��6*�N\�I����^���qc�t�{�k�y84����{_��R�41]���`~���M�L#wz]�+z�=�{n���������v[I�'�noM�s�(�z�p#�Ƹz������m#����FB�KA9%�15�1ME�X-���r�,Ւ�5ڛ���а�5��nP�	m�ګ���y�8�m���.v�yh}a�)��l
�+�b*-��δ������Z[;l��z��R<P ���B�]����.���l�N�q>=�������0�o��ϻ��no{w�7%*�>�����˶����Fc=��^�RV��(N4�k�yvti�5�պ��0{\��=�j���׷M�x�HR�k,�<�jW�B]bʗ��O
*Ƽ�N��ESs���k(�\9|���8f�6���#��^�I�ݗy��i��3='���<�+��ñBū�nIER$�y���"�̻��68�#�Gk�-o��g<��˯�q�>��|w!���ּ=��"/�_IC�]���Q�-�qcY��c2G��Z�{���z}PطZaey�ef��SW��u���%���/z�kr}�W�.�N���V�ߌx���BF���-Ϋ�һe��s��FV])�%R��:�l�.*ݟU V�PȂ�s��o�dN��[LNvgm���d��\�׶-��3�.�{H�ed����~E"T(p�n	8~�ۗ��E��r�Əeza:�V��g�M�|����s����`����~X��O���H0k�ˍi�xVDB?�+`�(��sW��.�w�%榯ǳ�y�t��~�ԃ�R�u�s��*����?�Ң�L�֨��9{k[�Gc� Ɖ(m2�)w��9�w��3zU�3Y��`����,�+����~�7������P��lp�B�o�BTbbS��msvu��%�=��ac5�j��x�)����x���j�`���eK��l^*�]y���ޡ��Y��������9y}Y��3�ǵ��fD4�]�uY��b9Gt^}� ~��/�R�v�{(w�-~E/P��4HC�T��:�U��̺�f<u��ks�.�45մ6�m�E�v\鍘��M�����b�=�pGۮ|�Fٔ��{}��+�q� ��/2j��&p�1�9��Z�X
[D [/�M]��	�>�����Z���*c5�k�7��0Z�7b�Oc޾k��:;���K�N�34#(��e�o�����6�Y+V[�Ϡp���ۮ��ƳC��c���"��}��j�=�M���y�~�᷷�!��lT%Ц��]ڰ��?f���_�k5,������Pz^�<p��l�~^<��3:���W>��s/!����Rc^r��=�{�s�W=�3���']q�@q��?����y��3@������~׹ST<����9İ�{�v��2z9��%WF�C�`j��	Y�����v,XT��ῶ
1��U4�[ܥ�8��cqb@`TqP������b��>� д�v/ovKB�!*��Q�۬�+# �l@��!+�r�0K2�6��u-v#�
:�����㌛.F�]���]��xnf`fhlKfn���n!��(=��oZ�]u��l�#��aH[�nݍ����%�ѥk)��� x��$ ۭ�-�f��msH�=��cZͲn��3
�,�^��[���:݈����7�ZVݶ�[�$��RR�[0�ƅ�.����qc�rX�[[$.B�B��)
�͔�Oc��t��$���e�j�j��T-�\�3-�e`R�d��~~�.צ}����7f^���/X��뷻b����}�#B�s��^ֶʟo�$b�Y�*PMDB���]��N�o�F�����fw���7= >yKU�a���u�����v��+����R�Bʃ�p�a��QB�U1p�Nn,؎gsU�ۇWY���۳U������(u��q���q�iok��x.�iT-���p�j�c%$X��Gơ���m�����p�dԻ��y�~6������e�e^P�cI�7"�`�Y�G=[!�iFT�P�H���Kl��Mn"�� 3;UjsަԮ����^�߰׽���x\�zE�=[V$�^�nP���M�s�~۴���S�]	��&]k�;i���R���*-�CnV}Y@>-Q���M�j���Oc�p�b���~-t�=/�xӬ��|}���K]��Ҵ����'<����v��le��Y%K���h�j�m�h�l!��4,��yj�64��������������4�H�O�ж;y��cM1-Z������r,���7�W����l����~�U)*	[���pܻ��������zl�^�����]	L�<�9�U���j��n)�-����U��0I��^�Y3�o%k��~��A����>�q�\L�9��.#�:g����m3�;c�}�.P�K6�ORά ��G<i��$
m���cI+7��N�x���V��d�s<�|�2�i5u�mn��l���^iǻL�4N[o�+ї�4󆸻����!8A[h�����_��w��V)���˃}������4K>^>�{��^���oN��:�u��z��WA�����d�1 �TQr��L�L�queo�ű�eDDvp�9��	t��䎍QH�Z��w[��{ǌ�9+3��g�g�X�5ҧ��EK�����1C4��O.�^�/���u���j�A�J�7����o��4�>ᣲ�3%��%-����~^��T�^��Uc7՘�V��Yx��T�̫V��v{`wwu`]�h�Wj�
u�{�3�c�¥hbY�Vk43�7%�b�YF��E����k���ugTŖ���a5�K{=
���Z������R����W�].�6>5v�A{���N�%!��ڈ�=���Mn��7f�.��wV1hL���HM6�9�u�<��%zA������nF��헀n#5x�����\��x���ʍ�}����g5��g��t�Յ@Lr� 4��������9���op��������k���lv[ٞCU��7�R���*��<r��;Rr�e�B��1#x1� ���X�a���\�ZJ��%!�6`��M-1	b]\�]VhB�Lݲ���&"�S:F�����:�v��F{�h�S;�X{NxwVK�9��]^jz�k�֯ �>�堚�x�ad���ak��sz�:���_�01������$��l��}Y^�����jm���4tkTqW���6��lӢR�*pCPZl����=�N���x��2�Y�^l����Sw��&��5�ǷAk��h��X;Q���xk,��}�	P`�4�)]۹���T��*��S�k/m�;��G�ʭ�d����3.�&7/|(-X*rn���Y":�L��/��3@Z[�4��.��e��S�ڱ���E��2�&��nƫ$�yj���m����k�����΋��f�ķn0�UL��@�� GJ�Yc[o�j,�w�F����W�t5�]��{�9�Vq�
�)�m\ꗣ�y�t�z>�ŞQE�(�K����t$�
}JLK�JnY���-��k,nr���li�Z��lC&�J�a'	��0O��&��ڗ��_���>�<�"��&n���>Oݵ�'+su�N�!cQ��A_�ji����M�o�vP5��F��t���j1�/�jtkF�g?^v.�۬��=�aW&�E�=�%4��ͤm�ظ�>���y�֌gZ�X���i�Z���
=}��
*�=z�<:=1Z��j�b����qre#{��������Ɗ�����zڝ�����{^e��!W)v�K���y�^\.��ٹ�"k���/�v�v�F���R���bvD�B���wi���q5�~~����x�T1��-���L):hm
9;ncf��͆~=.�Ӟ{:��ru�J�E!�f�s�R�m��A�UvOV�.��֦3S(\޽��eC�N�{W�\�+Qͬb�0l`�ܾ�koK��6__�����r:i���f�\<�� ;/m�w3b�9�$��od�Fhִ[�������o�e2��P���g��]l
F7Y�Mp�L�	YL�Y�6n�@�uav 	��.�a+/�1���4�n��vmR�n�THͶ�kz�@V��������B%��4����ɫ�0�aZ���xۈ!��1�+�pݍP��]s�%7`�j5YVИ��X�hB��4�Kf��+-�Mx�����[oim�v�1u�	��&+q�L�]����uښ�#o|)踬�|eb��"��;Ri]W��1F�$�R�;5�f��K�;�[��I�ݼ<��E5V�Oו
$B�Vns[���q�s����w�~w(	����Y�07�.�}��n��umn:�	�& C-���7'D]��ifD�S��ڵR����������A�q�%9�����|�`�}N{Q����,FS��'Wyh�33���P����L-loB)U�{B��r��E���~tEMZ���rb��o�;V��= h5N�u��K=�Q�N���@�
[I�S�\���=�-��۩f�3m�Nz������}�U�5�-�;�w�:�:{�#7��|ki�D湍&t��9j7��a��d�f�{џO��=������&��7|Z-�quZ#c��v�ڬ�fc���~݋��v�y2+�V�zd�Զ�h��G���PvK8s21+-�1[c1&�˶���E��iuh�Wmt,�
����_z�]*�5�%��q=c�ǆɍ���/uE��G�j|���ff<��a�g�[�W�]v�µ� ��7H;WV�6�3�1ۗ��hD���^�y��}�;
Y�&<�U3���:��f��*n��;���JgK��2�r���Ⱥ��U�5|`�m�9�]���c���;�{f�� �(��җ�K����}/�?OE�u�}���k����8;iiQEA��@1Y���v�:+}�3����ݹ�=NHd��Uҳ�:9�ϻ��Z�(i�of���K9�o�
�<��v�0�N-��S�ei���=g"�1���IN�x��#�g�	�������>U,�(D�>�La}~js�d����9r׽Y[F'���A�`5�w��]u��su�/;�]��%+X/6��_L3yx����t5p���+�&#�,�S;U�靰1�%d ��^]��~F{�0D��E�,��WL�/i�ufmG���m	l&�\�����f�]jBc[�ɽ�:��g5x(	�V�/z��C��[f�L��$Y��}&��u�kLD¼��)�ݧ)�`��#�q����M �h��n�J�[U�6v���o���]�nL`�1k�M����"+���6��Z��fT콐sW���[�3 �N�]��ػ?]�SGR�QmA�E]���)Vp�w;�=W{��m��ĕa��?�v#���-~1p�����}M�ْ��QĲ��b5�9��N��b��hD�u���c�.�Sn^Yn
�sm�L���y.�^:ڟ��[������-��םS��sM�@�Q���[8oئ��e�J9$��<��*�N�'*��w��hɷ�gr�q;NZV��j�Cu2�1���oU!���o:*=r��"�g]7}�|ޫ ؕ/�j��,�������f�ѐ��0v�5����t,���b�Gm63%�]���P�;���}׹��i���hN��᰺�6�n�����bN�*6�������vFΫ.,;��4��45#�,̷GDUɲ��@��N��v�7����-ܺ}������y������&3���W<ؗo(fqי�\�n�.<���w���GRz$U��_4�T���+0�M��ݕl#S4���/d���_+���ƭ�ww]��"/4|u�]�Љ�v��Yx���\S	Tf"��5�9ҏY�[��+B���%��hW�5���r�y*֨qR�.���uՖ�����0�xUj�wX��_=�6�q�$����kʑ󣸍�v�(���pgLU�u����4P�/�^��[w%�ʚ�w���N��a�ܷܕ�QLneuMT�w�6�3ۙz&H��B��L�͝��;xM���wyۏW�O(�K���2eݕ4)�̋)��n�s���$oYɫnj$���Q�2�v���y�<�۽[�ɼ�H�fL�(�!���Ħ���Y�^�M+�i��b�����*H� �v�(#��*EC1QwDS菰G��u��D��g��u�rfU-9�/���&��.��Y��m�DC,��b.ըA�U���'zDi�a�sc$�~x�y7ݷ�g�6��6 ��5@}�D-�Q��>'R5��z�ǥ�z��"����g:��}JeZ��P�J��rg��^z��ݞǑwP@K�8v�}��{_R��h�r��(�u���(��9۳vj<�Y�U x͑���h��Öo��dOȒ��֦X4���s[omY�
����]�:Zҙ�@�l�Be�c���=k7��=3�=.�xX�@��(�uc���2���wm������n�ﳤ��Ӊ����S���0�}�]�rl�
�Y��0��2�j2� F�����*��`���L��`ͮK�wx�h(i5~����lC�=�ߪ����X��罠�l���Bh
be���#�޸�"~`6D7EK�;��>'e(�����#��Y��(����_h���~���w�㣐A�ʗ��]�PX�wX��]&x1OSӊ���3�D�n�7Jeɚ�iaE��޹��棼���������L�S�P��+Sϲ��3m�\�Zd��~�s����ɩ�U���}���
ͧ��ɮ��2�
j0Vzփ��Q`�+�K������K��U�����Ȝ )�����i*��̢��Cb�G��u"��n_zo�{�F�i&�%�`���8t��9]��Y�q5�v#��\��<�9O�e���f�*��}l-`�=M������M �Ϳ �'!�@�z}����rP��\h�WCP�5���f&��Q,ױ�f�D笇["���P$�#�,�{ϒm��x��{ʩ�\�7��4�y[�l�p����U�8#��n��v7=�`C��*�L�H���'�Qۈ���C��D��Q7iJ�E.�αy;�`̼���y}�F��Y;�6<nL^�]<�>��'d�nB����}�⽧�
<�C��<�JQ�0N��}�Cx8�<�8�@N$
���c� �&4�����O��}J.c�h53���Ez��y"�ֆ7�0��_;��w�aס�F��v_yן.pm}���.`z<CDCL�L6ۉ���<�NXz3��-�g����F����pZ�ݯh�C�ո��{k�g�Lf�Þ2-ߩ�uvl��M�����(�KT�	Y��K�XE�a&�MV�-E���_GWb�c����-����9��3�&��:5Q��
6G���fW�J���0��XpbB��Y��|�?r�b�o��3/$6�Ъj�߼����!���8�����Vf�̓leb�[H��:��A�/\�I�����)�7�ɘcs���R�0l>bm�l!�Tڮ̋wYm�چ�Zc���f�dn��B�-`�fI��Sz�������jZ�Z&7�iKV�,ΊP]uWp��m�RіX�1Jڭ������De䄱��j[] �����.�5��|k\�T�pY��n�v543M*�����˳��]Z����T�ͷjm+r;1[&�j�Ń�7WM)�1i4@��Kl�
�����,
�ˠSA����,�pxń��6{J��6��JLme��32�e�
�+-m@��[m߿Mr������ǋ�m�\����,�I��|��Et?��fI}�Z�����κK���=�ed���O{���!:K�[�p�#�-c�u�2�y��93�����ڧ:���^ ��`˼�5�bDo�g�yo�׫1�zN�ܰ�����O��I�oЫ��p"M����0������۾]yǱ?LD�_Z��ǆ��ޣ�ܫ\fVz��k~=��p��y������
�����1�������Y"���'K�Vp�>yz�Փ�W�'z�~�n���|�3{r#Ӻ������ϧ�Y�2�x�Ðȉ�����A�|e��gR��ڤ�Z~��eCb
�e>����S�d�V�*\��L52c��zs�eκ�R��GUzH���޳W|��؛`a��R��y�W���}�n�u�:s^�w�:5��"�qJG�F�dЈ���̺����kz�
us��n#.�rYv�e�BLH�6e��;����aX^�`��ֽb�����/�T���X�
��S־�WQ8�=�C��;��ڼ�x�d\gFZ#�(��N �%0�� ����9�����i�^x���$������v�\c&mL0�m�W�8�{��xi�sp�l��U�J�7��Kǎ��<N��l~y�M�tu�cK��f��:}�r0�M��!uWTȿ�,T���X�WtNv`ϼ���&+Z~������)��W�(8��^D�y�ye����4f'	�T��n]��q�D��k}�X3�^��#,���w|�]���J���a�_[��S~��r9ή�W��vKY  ��ŌY�=Ѓ�{���t�f�,�=;��,-)ك���
���s�J�i�1�ܶ�Եu�V�w�5wg���\�r�����D���d����N쩣����9C�狶u�;N����{֟dv���+��T�^��r=j�kC�~u#��I8%�u.������J��|�p��Ä���e2\���m���3)f�,��fgLᡋ�v������ ?y�j��E���Q�Y�CA���{��w���+.K�z�wc��i�Iʨ�ˇB�PE^x�:��T��o�$�3} ���h�LѮ��<�{eX�����9��}��$v�yLU�\����0:r�Ϡ\�U�8)3]n��S��~������;�aL� �Er��l�F����8��>�T�/3�Ov�7:��igp�_k��65��<=�>+p��1�X�C0Aze��5�в{��؍�ϖ>n��������(,���ls�u tc�-�]e��fǛF�(D ��~#���Nw���0V{�BDv{<��������̅��nP`4��IԌ�M%3|w&���c��hM/�.hǉq�[���_�Mt�Y;��g뿴t�XB�d|#-��GԻ:������){bV�}���x;e�
�+ �ӘS�����0m4~����/��C� �3>���<���ꢫ�9cn��=�"�ɰ���z{�M���SG6�����ZYx�B�p�	����8B��Ѷ�dve�ncL�6m��Y�3	MV6�m,A�B֫s��Nw@�^� �ܘ^��|7�[��P)^�"I�1̈Wn����ul@��6��\!��8������]?���\綦�e�Q�� ��&�tw���{3�}��}X�(��1;�֥4av��*��!ٌ->쨐�:��}e`����÷׊,��B��߭�Qʹ~��P�G��(�CMՎ:�+=�xQ��u��D��dO/�_�:�rŽ0�}��vͦ+N�Km*��F�u�a�;1�l��2.�1���z�
갖�
�$�֊��<���"��3:x���-��H5~WPj5���[�@vd�`=�|�/hu������jz4�o�ш�fc]Y%�6m*Em�.mߟ�X�AGK��%A蕽��|n���Nw.�̲�*c����}$;;���n�:��d���u̾=��F���v_:���h�5�'��9S��wt��SF]��y�7R{�z�W����bŒǔb+Ɏ�<'<C�}3]����c�*@���NǷ�_v�?qҽ}n�-���Z�R�!omQ�U�l�M�d&�K��Fh-Sjl�e���D�I�#>���*ͩ�y�vI9���k��A�^�͚gf��{Ňؠ_��.�Q�1�o��<`�,}�[[k�����(z)x���E�T_�	M��zO)F��">�}k����#�푩�WH��ډ�.�>�����(ݷƳ�G(���}��ƅy��_�u�k��F�� jBjL��Ui6���U��F6W[�����/�eɋ�Q�y�b��B�@!�1���V�3~�i�	of�\{1v�lƻ�@�O�[��r�|�H�<�[0 �NEÂSq:.���wwu��� �'���n��*��խ����n��x_U���:e}�E�ӟO,�kdMo����ă[����{9(���v�+������ead�X�쑗U[>�0kf��s��#�co	B��,G��^t�f[��qW���d���)͈i}��Ko�i.4��j�m&�Zs��e�0��ڐ3㋺���)%���z�}�������[ڌ�k%L���v�M�U��L�s�r�.�yOk[�yQ�9�g敚x�L}K�g�ݻ����Hr��><��(~�bb�Յ(�@��Yql),u�L��lUmΡnʶj����7:݇,@�\Y�ͭ�l9]\:f��!n��Ͱ�ܭ�<��\u�;K���YVX��˳��M�J[G\�L�R�xDX����1��r��-�u]-�41�`ue*���^t�:X�cl�]�6)t,��%Hu�͈�,�-C�c�٘��� `��� Y�vı�&�ۮV�͛X��1�X���ɥ%���Fٴ���aB���ѫE�\6�v�UNRDU?���<^I�4����7��2���͘p|������4��1vB���3�<#����qd�q�^���x��B'��g3$vmd,��["a�%�����Zl����t����|gO{L�_ݽ|R\S���h=_M�'�����w|��/��%t���y����q�kFo�n��=�j�A �2�m�����h����!^#)z���M}1B�i������O(͋*o��޿&��n�k���������,�|Źc��	��8�ZMI*S>���m3?V�Z���:V8cfa�'���������g����B(w�d'�25�k�~Y�5|xt�U{׊�=�}Y=1�μ
yݣ�S�ߜ����+�j:�s���sd�ly�o�s�X+n|�o�8��9\�UKs��Ks���sq��d�t��_��&��QZ�'睷��e��g��q^��#�h�Ӽ,�&�j���[K�v&q1�����F[ʻ:�z�b����Qj�&�j@u�FR���dd��=�O��݌��p =���{^	���s�^͘�'b���ߘ�s�$/����",w��>�9�|Yim���2������]4��Dwa�B+������Iu��y������Y�ۜ �X���ef�ۚghyY2�9Y���uc���v:`���el��嚙C��f���.R���{U٪���ͮ�UڔZד�^���Wc��&=]q�2�=�{$n�s?'/�"uR�J��dQ��r���v\b>��"��jS���M{��*�-��<��77L�_�)���ܥ4��EX�Fs'I�5άz�a�M&m���J^{�vw�{]� {�5�m��V�+�����{k(���Dw����M�_���UJ��� �3����yl���Z����ɘ8%ast�kؼ���'%���him���MG����v�P�L�+��;:�*�������4L̙ۥ
<��u:��5P��G�)�������슱�q���SDݎ���F����}��l̥��g4�T��ky�k
u�l:�K-�P�2�[���6�i�L�ov,���FU�H�
��8��hY!�SV7�U�x�0�*�[��w޿n1��v��r�Q��6�w_���(^I�F�"�=���5F���GB-m�X7R��F9�����Σ�
�}������9"��2�u��b0#	�񬐍��NNAQ.lx�ewϮ;�p�vȯ2�P��N��\\��x�#��S��>�ޗ��֡|0�]�z�o�dY�ټr�8Ci*���f�M�i��HZ֫�^b���B,�1��6�D�����"[�n����j�jhҮ����R���x-����o���v/�쿣���+��������޳��uY�H��"u�"���s~�b4��ot�z\H�r�u�6��r�"�"��	89�+��:�ԠI��^�{/�*�ϢR�Х4cԳ~�k�{��_W�P�c�_,8�A���?"P�2Jq^�+j܌�6��/7W.=�	�*��C겇)�p�q�+��bL�&Y'k��Ww��,�D���<��f���K�`F[���cM�jR�͕7�'�6�f�Pڴ����;M���3����K�bm��cK4,��Y���iu%��E��i����"b��*�K�I�l��LǑUk{��D�* �K+{�o���q�u8}Cds>�,{}\g�x2k��Ѧ6�O9@�eb��;˿��X},��9U�槔�Q�B6+���u_G����[Su��-��X~����a�>��N�u��Q4FL��E)�]��T�[���9YiI
B1�<w�oe�R�2{�]���:v����i����Uf	H���x�����Ʊ�{c���� p!�<��������k�،&�6���*F�>������7��!m�'Հ}��I��;�U]Av�z�>q������j鎿V9��ֈ�3�f�F1�~yR�!����\CSV��d¯��VŖM�O^u�#��;E�,�mgE�Y��N�o����P�ڱ]#�N
���{Sd������&�9yV����|�"��Q2ѺJ Li5��RGM'�c7�GI�;�;X����-�o�fA�G�Y�8Vg�����DX�����yVW��,^c^���ֱw���-���X�G�V��)�[��!H�Rݶ�З^6��V�:�j�����jPNP��� ��o�V��f\�_������(�{+���w��]��e�b<T��ޠ&��蕼"���{ ��g�θ֤�}���O�!޹n�ˁ���[�D@��9܌�z��q��c���XG{2`f}�#|\`"76�:�P�F=�}mh�_8�a����"b�콋��=7�u�~{$]�>5D�����]�!@-0[U�����$w�����2�^��.X�)��/�Vq9<ǔf�x�gԽ�<J��`��Da9wl=�x��~��lY�3�zmxe-�Q����Wz�*��/r���;�T0����%g�����s˄����71���|B>:��A���j���tv^��#��"~�!B
����d�� l��۪F##�O;�Bm&�=V���x*�#��[0c@5�sv&��{ ���&�
�c���jk��I�� ��X��� 	>����f�]2�����Y��(z]�Y2�+j^C�͖�j�y{����0�nZ�+{��6�#��,��m��z˝];�᪶�Fp��|�Z���Z?��-�q��}՟���X�\q�YX*&��jf̲j��ډ;��i�r���m��U��gw~�s��4f���v_�ʽ���zgg幛�sƯ���=��%��.[��gb�Vk�ِ-��We��j:ۅ�V��Y4�F-�;jl�C��Y���&B�����Y؋�D��� 8M	k&��慊�N�� 6,7e���|)f��N���� �Y�:>ss�A���v�b��c�{D�|��6>����R�htdl�~�	;F5z�p�^m��G+J�~�ڦ��\vVq�r�e�1��1P�9����4.��ܩ�L�	b�����ܼ�;'�{����t�爋�^��"�Z��y���kn�s<0��S�l���7ltq��v�m^j�8].N��\�藗sw�Rg�qm_�&�Kf^zS1�R�P�֦���\p��������o�wR�c�k��
���Bŗ��8H�]1�9\B�su�b^�7���P6H��.ټ͵�;q�㙜lhoL��\���r���٫Tcs�[�3���V+r^Ȅչb'P7fu���~On�� ���
÷HAL�[8
�r�٦-RN2 p�M0��%m��=3�d��, ��⫬ep���;k0�|���W�cOfU۱�s{t�Q��\9�3O!M�,�ާGǆ���8��K8[}k�y�
���DrHT;P6�\"YM��*���-�Q�P�P�i0@����0�Z�bK&�/&WTCZڻ[���%V�XL6W:�n��]5vWYZ3b7Yu�:ݐ`)t�����aeD²(墖j⦶��9�v�����]��킵�e�IHM��l��hF�e�m�����vQ6-�Օ�pCh�#���Ұ
�H�1�H:�u�f�]
gf%�ᵛX"�BkwR�d�-�hs��[�e���j1*��d��VX�:֍��H6�к�m��l���fݮ	j�b5ୗQ96nXJ(ѷI�n��a�l�֦Ű���W[�v���9�LglDm������bbk��k^:���M6�ٯf���h��jX<ƣ��S1����1��K�c�	m�Ŗ����:��{H�AЮc��1�� 2�!�vCc6�Y�X�v�)�[��3�54�(Y��:�T&�L�]�66P]��ZiX�rHº����l��u���a\(��v�V�ծefk����])�HU5�GKf���Kv5k�sv��բXm��4�5����p덥�^���CR����l������k��Ma	���=����D��o]��fi��(�S2�vD�\!�JK�V:ilk��	c����3�Pu�Sm���mYIL�R����-���+j�u����a.�7�zX�_3an���d��SeS]Kf��דbS7=��Q��H�i�[Y�iYHh[I���"Q�����o&�-u�.D�Y�n#���j9��M�K6^v�mIe�B�h��mݶ��Ԣ��=��y��P��l�M�[!����m�.�m���),�-�m��5�v+R�	3�ֶ�a�k��B��5q���M�Z>v�[��#�b���ŗ�3��-q�nuΌ)m�fZ��ڧb����lj�j�*M*Z��ԅ�CR$��vaK����Yf�\�S5,6�l��[�\�&�)Z;J��A�!�ۭ2��v�-m�Ѷ����:�f0���j5��9ܮ��j�%v�\�[L�6S3��J��n��(���L\#A\k���	�J�Z��z��^X��)�D�GX
�"`�#�*#� ��A
�ӺpI'@�$��}8�I��&�Rak�-�Ԯ�6��۔�h8i6kn&���MB�(h�����cIm���_���V����l��Cb:i�^Mu���6b��6�["%�e�ˮ��n��.��je��Z��d�S�[R���SSMZe�x�5x-�S	t��\%��˃��CCL	+f��2��i�y;j:�����[	\ǃZ6���\�l�2�[�a5e&��)�tY6�����<�@/-��c��-5+
M�9iՅv����b��@�.�x��Z��R�h�R����nD�*���	�����d�g<?����e�oy~Lw^]ɛ[��|�3�y���V�=AH&ۂ<��b�;�a�>����oz���0,UIc�����ok�]���'8�^{��y@D���,n���G���)�Z��y����<���>���&�iq�}�������E���VzH�%T�2����+��l�6E�{�X˄1�"I�����uB�Ӡcvf��v|E3՝�;��TxY���VtUaJ���7�>�p+����pf^_��#ᵟ{��ʶ��3=�z��Z5�n{&�>4����{%��R��I6>�A�s�0�^�ۋE����mŞݓ�W���FO^kdɃ��ٯ��"�v�(BQOo����2c�4�x.�T3�\ !�k':�ꎡ^O����n�P}�<�P�w�P
�W�_��k��i��.T^cL��C���{�����4�"������c,�;8��mq�������Yy�bl۬۴#[�^�m��][�A��-1�����UP�Y3����Ƙ4{[`�7|N �渇|���i*�xS>DGwj�;|3;��^'��W���\U=B��@�����x��0����+W��6p���	Xh	yCY[}n��povm��$_A��[����lUV2��ӻ��� ����6���_��Α��Gil��'�Q�2�y�DЋ�H�~�t�������cS[L��Dƾ���5M�^�Y�Ym��W��j�ꑊ}�K��:BgOݻn7uA?�����l7v�����9��֧2nY����=��˲b�3�S��%Uc6��Q�v�3+�>�W3*�蟚E�!�XD4�"�y���b�g�7��ҏ��^��N^`����h0
Q~���:T ~����:�<��RGI�gߙb��A{�����a�l��͐G|�;+�v�qB����_m�7��vK��t�^R���P%[�Ak)�qAqV|�}OޟTTU�4�[���޻X/G�)EkS+e��^���F�UMt��Wm���Z�vvc�J#�uͺ9��V!e4n�ge�i�*M.�m�5lmt��HOW�?hhЃ=��b�!M܅'�U������s/vk�A|q��H�~�4O#�;��0ֹ�1� �j*l
i7�P�Я��3\#Y��+:�{��{QP78�]�X	Q�g҃��� ę��F6�u����\���ƯuO�o�����hؐm��p��y����s\ds�s՞�Y�8#`\ї����/ ����ɜ�`�G���9[����ts7�74w�8�7��\'^en�5m��y�\u���T7kZ>��b߲�{�j�; �L ��a�NMt��U�ז��׍'OƢ%�/�A����7�Z=%#�A�^��H>&��,���4_�m�Z��{}��c��lY�,ޛ�	�`�s�{�O	���E��O�C0FZA�]�j7n)����s�Ú���~�o}q?L!��	�YU�]awc��ݬ3@�Dا��p#�W��^��3��w�.e���xm7�@�%�������5V�n,&[(�.�64�m�cmM����I��&�ݻX�X�4��ڍ��m����81 ���ARL�^́
{��oq!�MΜ�;U����S�ԁI��D�2MW��'<�~����nFf #��4 i8I?�:L!���/㴇.UUZR�}��F:曗��Ig�G����s��[vf�JhZ�4� f�PO)�2*��m���m����u�+ R�zK��2��r���g��N�J��~��#�Y�sL��!�|�>�?v)w|F\0�%��f�o���_"'1�C���@�q5�DJ:Q���Ln��i8M��\�<޺�
�{���.����eW��A]�-7QUw��:M�v����ʻ�#�vo'�
�,_*�N�����|t�"[� �{n�i�84�/6��Iu�ǃ9S�:��0VO;�b���=��>����a��%�H�:S	wK����G&ns���Wy��Pp �$+�����w�;��͗Y,E��Kqޮ𪾤���#	w�f�*z�{����R3V��{��3YU7��O����]��\�sb�hA��J�W]��6D�ٖf�Q��A�.���SJ�K�m��ޗ��wf�\�׹�x��p]󺳵9�֧ٲ[��H��Q��UG>�!F���3���/��5&�;NQ;��\Mx:Ů�<�M��#�)��J�^�tyBZ��(�_�^�ۖ����;^w)jY��5g9*�&�͹�.1�j��Z'�T^��ث��-jj��������B� ��n,q�m�~'�&.dY3Yӯ�ǣ2[[��,(�4Iu�.���r�ߢ�޼�w�U����Щ����R�34�ޑ���"�׳�&�hX�	�(�Nn�w�];��B��<��ǽM6?k~ϸ�~�C#���^�5�0Y���R=���[���fs����=��V���{�~�jT���_-�R��	�P�Z�r��Y�17'ܷ�o���Cx�dg]��^h���� �}﷯$'�p���f٧��m짫�Qę��xV�0���K�:;1^C�A���Ơ7�#���a�̩��,Y��Ov��˘�:��M�����ɵ����t��Q��K�*�k������$��9A!$�lخ��n�5��V٦J��!�q]���Kf�����k�)��^��u�De�t(hJ6�������ef�@��V���L79��+��y	eΪ2�4�KKI0�&5��V�Z^ٛi���#��\�t�u�)JPh�:�F$kM�KUƆ���RifI�6�њ�,bL�fڑ5fvK`l�n�X��f[�ӫj��.�V�%f���>־�s.��R�k	�4�ֱ��H7S�����ƅ@ݢV�քx[�Κc)n�m5qv�~�;�2�������ʟd�l�>�ɫq�F�ũ������W�U]yQ�pu����a���ޭ�t�,鈼y��p>��@8!Y)�؟����9���7�.�s��[Oӡ��?���6>�J<NFR�v�z�њ�  �m�˨��b��XuwY=�+WWw�!
�Z��Y�������*��lϣ�M�K"������R�>[�P�<���D�3zch#��MT�!���ngO������E]��6$���2ۜ7J�zG�A|�ּ�b�p7*A��b�t͓��t=�n7Z�Pk�r�K�pG^��Ng��8v�_�����U����S0 j�]�� � 
��,2����grlj�m���{�qX�mxO�%���ջ�3s�=�fF6t���|��l/P�Ǖh�c��s��ж���~;�ݩ�Xk��Z��_��C�N;F�I]5�.�-�軲���	���W���]��!J�c�( �E��J�1e
[�å�X�B�+e�@��#�4�|(���q��ǖ��sS*�o"t�����C̻H@m#c�P��$j-|���0Y)�
n���r/����L�a$�u����	���
�E鎨��gJ7ݚ��z�]�ep��k�s�B'�)oU��o9�d؍Ư^.�{������,J��&�s|7l���e��W�����J�S�o�6��j��2^\�t��h�q>B0�~Z=׎=\V���0�q���E{�/�ncns�M��d4�mڸ�S?p�%��ݏ�='B�Z��c2{.�����i_s��US_Z�+;%���!h�31����GO����&��5�~���=;/� �d�8U
�����Y�뗮p\z�z�jz��H��K\h��G��p��0~lV��̋h��Mu�1{����-��U���t�;4e��ذ-z�� ;IGb��v��-�_?;txu̱��@�͍>�e��Xꏣ�^�����~�^$@���z��pU�=�_uW뜥�\^���BH@���a�n����W]"	��v��mņژw$�5�����/���1�";�c�ͭ���v�r��Sw��K���<k��Vu9�21�J.�r��J�癴O��d��zⅈ"!� ����c��<o7��C'��d�Zp�-�wdѰ��6:g��Ðb�&�e���q��*�Gz|�w����2`�Kb)��@��N�;%��r{ƻZ��3�<�ck"�t}&�Qя��)��i��Ԫ��@�}��=�U�?�E��~�x�Xo��@�P��B��y��/�]͂ɖ"�7E
:���o/�Qe��ݞ�$���Nڕ�]�LO5�U�u�R��ʛY��37&$g`�k��B�J[8ݶ۾����Vx����٦����m����i^p�F��d�;����E�E>JR��o1���>Ύ�����E��6M�\�m���g)��	�N�S�f�>�f��%����j�<gٙ��ܗ�qq��w����Y[B�Zo�jnΘ�-�0n�+��{/�B�E��C�z/���qW�j,胔���V���V�|���w9�۹��8`�Rp}�6ʊ!.���'W�V�Y-)k���:�c�ڗ7+�VWh[u�h\�n�Cu��m��CM�7d$р�d�l�ł�-	��zY�^�h޹u�:�E��fZ�"(�	QX��O�x�wg:�J��{չ�	�$|�*s"�"N
��~��ckc��������5]˝�y��yq���{^��"��L� �p�}�{���W�4V��[��i�y��c�
<����}��棉���\c���!��ue�<������±6�ƭ��6ɉ��v{ɏ���j2ڵ��H�@�����X<8>�O�e��i���N���_9�>_uM��4t�
�5��5G����Z��[���c%+QЦ�w�..5���ϳ��=��3�EҬ����))��8�X#��:��u��$4M��
�v-�g�����_�^��Ὣj��\
����2**����_o!�t4�m=y���ڒ�w��VQ��� 9C8C�u}u����WԊ���;����>�T����}p=�
p�Am���mg����uR����W�����G�oW�]TuQ�+�3��5��^~}1��)�^���K�U��k��-5���*��=滚�ͯ�:���є5��lG]���e&�.u�ۍ0f/gH�(�K]��VGR� w���'΄lIW��t8ǨAh:���,�x�A=��8��G���&*�Ff���|���td�𱌈��k�{��������E;���e���m폲�3�ϫ˪<;�ޱ+]3��� ��h�Hū)|����*�3\���=S^g�}�ڢ�R����~���t���;�4�YBa�рKn�q��I�J^~��U��s�08�_Y����#�qٰow״o���^����+��EV�#6�e�����A��V.�B���&��DS�F���K8Y�~�~s:�\_��u��]jB'ï���{�A����=��揲B�D�*�����I�`�8���%�J(�rϽ����"�Yl��yc���T���{�xڨdM�3"kj��s�̂Vh��w�W}�J�!��H+}=�U6��y���7����>r�������7���M|U���T��/�mlSٛ��f����,_z�5�!S��~��̟��V�x�Vq����k6�5�,WD��8�ܮqM�]<�[���j���F4�P�Y���xo�k�%\.�{@�H�VA���l�T�#m��.�m�P��h�ك�.�m��i����x�9)�c��k�Մ&��k��`u�nR杭27'Rе�F�mr�\2�1�k�M����.5*��6]��e�ˮ��f��6۫�im�n����-�j��f�76Sh+h�Z��̩y�1qR�T���c��k�x��\���J��-�1�Q�Mn����<Mo%mڙ�6�M@�l[1�|0y}}�*ӁR*:[e� ���\\����%e(���߬���lA����뺷n�})�}ڎ.�5���u�_v^��:؄ �LQf��nG<h.<��V�H��ht�eǇVK��i)�S��s���ݍr��Y��{7�| ���}7�Ϊ�:WfD��voxR�(�,�M�.���Ӱ''��>�U-���Y�l��F��{�H����L�����5u�i���'����t�ld���B�J{}Rꏒ��0��dk�p[�n�6GJχ�3}��+r��ߍ,�e�귘���ތxs��(Y�Ueo\�e�>�&H���貳ˊʇ6*
�)�+�X�x�us���;4Ϩ���+�s�5��dK�&�M��b�����hV��dUƏn]u�˫��D5)�G%C���?x�������7��ύ�)W�p����/sF�g9�d�>�nv�ԭ��"���(T�^����+G)�	�dm^��J���5�C	�p2ܺ�)XZQ).��M�eln���X�)n�q�V�UJ�1��[E\�)9�طv��`@��6��h���4�����d���|a��j޾�nG��cS�M{���Ф�z�c$���4-�θ�Q�σP�E2
����3S�Y���Tv���y��s5d�l�=�t�N��$uԌݲ�k���@ul�ڭ.�Zx���0&���ދ"�f��������u<�=�w���i|\橓�=�륦�;ɾߔO׆� Ӑ`	ޞu�a�[�ϻ�Lު�qg��鷳]~�3i5�W�1�(2IGJRk}y�
7��r�̾��e�*��o'z��N����7�kǮ(9������t��+U����u�{��0+�Q�z���[�Ìdd�h���,�v�<���c�w�dMr�Q�����Q��W(���u{���^rɲ�ӪP�E�9�r�o���yU1�
�|9h]����0؄�0ᢊu7���hLt/E�;&��u�J$G���+1�w�FF�fᛏr$,J��w���XU�ح}�_z!\��jT"����lf�A�@T  �h�a��\��B���Wd�G.�1�٬�i�9�)�s�k��ܿ
�������k���~5�d�`xEoQ��g�<����j�Y���u=�6F}�'J��:���"��xGS�s����SR�(Y\��DJZ󘑾�Pg m�L��w�lnH��Y�O;���{ƨK�윃Ȉ�y9�k��+܀X���ު�מ0I��ȭ��#�W�.%�%P���p��r�3^�G3tN��������&3��k���%鸈vo�mq��9%��>
�W^p�A�3�e��l��1"��X���j���ݙȨmt��z���@~��3��z6�a�����ś˳,fV7E,r��f詝���L�4��vc�����,˩z,Q�ҟgT�R��%���M��ڼ��،��'[w�ʞ�<.(�ni�mFJ~p�P�X�����`�<S�Eu���Gx�v�g]��"e�i����`�;;a!��'�,�6��'7���e�p-7�GM;�bw'"�9�y�ɻ3(`����:%�k%�ه6�[� Z��gU+��IWni�Ej���]�����,�;����Գ��D����a;�O�()��],�9]$[�.�.�<��:�ё���u�S{S�D'���uqL3��h���*�i��Q�2�����~8Si��װ~U]��Y3�z�_w�6��oz��։#�{�����lg/��v�B�]�3;�"���uZ`��λs.]�����QJ�R.D�M��c-�6�{J2?��{�Q���N��qV+��Trꉜ�.��;s�V�U����X���Ǧƛ'�b��qj�8����^�-5׽3�n�k	�ƻ���¦��C;b�c���(SP���$���i��X���q�A�SP칒����p5���r���5�(��\:�(���Q_;�����֬V4�ֵ݂��;3]u\�r��Z[�ܲ��[k�R5�<���vN��{m�'M�u���b���#���,��s�
NY�V����G2�u����ٗ*�i1�E7AA\�� �*�CDG	���4�z��7$��+�L����Y�/�բ�j�zz֏)��B$L [x��)٨1;儙����'n��E� �%%�}J|������au�fs��G*�>���t�V˽����q���9,��~�p���$%i���n�3����o:�eU���E�y`���_WER��\b:�=c���ơY�c���4����1]��G氓�{q9(H�����E�I AG��ٱ�V�̱MRل�.K��Al4e����i��s��@�RU!
��P��}|c�{{�X�ǳ�u�e%�>v����Eze�fۄ1�{����F'2��PwpD�oFg��=�������U2l�mE}w=�+��(��o�����O�26'�IgD�D�S˴��5�m�ԗ{o�x_�/��0N�t��j�]��oB.E�S��c:ٝ/k��H4��7�*f~�J��L�C}}c�^>�or���H�Vy�L�Xk/~\}o]voq��G6̉�$�t%h�u�
�z�W\�6!�F��`�����[��N=�d���t�7�k٦��U��Dt��T�+��
%�:�6g�`_[P��[�c��yO{/���Ne��`��^C�sQ�.���tUi������g0m՗g����NGfY��	NY�<H���h	|,���g�Gڶ���ME)�<W���n
m�L�lMa5i�^L��EW�1��oR��c��oҥ)�����<X>~�s4�n�,aUmL ��u��Y$���8:|1����я"�����Lیi���b�'Z����۬�6l���ð���+C�3�!+(���uҤr/�)�2)vl����k�+'�K�ׇ�"x�P}"�OĖ�1���:{�W/Ј0mʏYk~�?Έ>�n��
ۺ�L���ܒ:�0(@	��5uor?�;=���]���f)ln�־g|�����q��T��ܪ�gY�vL����μ�=\{n^a�}פ�\� ���!(%�S�C%8��7����`[��5��;�1���u�b	���W���_��W%��Th$�c��k��e��!|��^�Z~>�;���&1B(Lw������t�����s��ߧ�� 9�j豛�e|#ϲG��61K�״$>��!�wxnc����-8j���`T|3�{uY���u�H�P� =}��?�/`�.:��zk�U7P{C��Ƕq������C�צt�Tؚ�g93��x� �L����-�\.3#v3;Y,�ڹ��s�,_f�gH���F�f�3*7]��iލ%�W�]/����V tA�1
ض�����
g9��������,�.��M�,�+W58�氓c1����@0̏�x������^ҝ
XV��jf��n��ń�B�ZaffA�1��cV�F���.�l�V�B�	�LXQ��Za�v:�e��V�<�b�jRTF�+kqrM7 	�a�j�D�	��#m5���Z�4
�����:�-�dշa��J��vZˤ�L�*k���.)�*F��.h�2�%���Xzn�:,�*��\B�� ۹��1L����ʗLKu4�U�	�@�IK(�A�7H���r~�ƾ��-.ޕ��5~��.�+�ߞ�c[����o
�ݽu�V��T�Eҵ*P◓��5�<���i���1�7�\�L��p�i���V�g0�ov������-%���%��ܨ�Ξ�~�'���	=�[ɱg}3��x8�h8}^�<+�҆mǣv'�Y���:��e`UQ]�e���j��L]�zǷ�y��Ĥ ��K��׽��Ӯ�����=�F-����^�	٭'���3Nu�VG���5��T�>>��[@U��_;8z�lm2[�3���W�ފ%c�w|%ذ=޳7��>�Q F�QU׆k�y9��x�@វ�;g[����^Ӊ�>vАe�G�<:-pTR�ZWV��$k��.*SZ�sZio?rU�q�+@��r\ǆ�`�.�+���싚������k���|���a�vp:f
0'=W� �q{�Ǧ��>rYe��b7뺜!�JAf�&K5�d�vk����v 5h �!2��U5(�Lh����G�&q�H�3o��W)��Lt8>33���
���[���}8{p��w�цd�V�ܠEP�s:��h\�%��k���}��i�
�6[sB�h�4��\��ʪx�"5��1���g��U4-Y����[�t�;ܕXoE� e���}BX���1���J|���z-�*�t�MFg����:8,��� ]�|pt!�M{՝.���E�$����ǂή�WU���t�O �ob��;;8��Z
�+,[�h�����~�u���yP,��:�dv9 ��5bp��G�_j*�h�>�����I�>s������U���J���)�%31��*Sv �숇� �ܓ��{�5�j��?kk}�Nhi4Q��JX�C���e)�������{4+s��7�ׯ*u�B�mIoأ��)���I�~�~��1 ׮��S�p%��<�N���)�Ew��|g��)�?LZ�\����W���w&!G��:�}Q9�}�wpޕ��(�YB�-�C��./f�u1a�5D��5��hs�u.�XF�ѵ�&b�	 M��0q�.Y���c�<VZMv��W\þ��^�nT��uU�mJ�I�>����≌�	jݼ�7�<�A���]��p�n`����)�1�k8ؗ��u�1T�}>�����&�ӗ�_̴�B]���·���f�
=�vN9O�u¸E���{ˍ-U��Z蘯r@r��A��6����[�]���jDYSU`�[h�}w/�yˮ['�t�sэ̥��2�}V�o<|<���\5e�T��V�8�7IKwMd���Ǝ��,�%K��n�!�����,@�E���tZ.�t�ԝ��E����8��~��2��������̉L�Ŵ\�feBP�I��l2lw�J��:�Ly��A���<�|c:���؊�Ȼ��M�v���
{��.{ �ۻ�؊�=��b�{[ ��-׀g��5U�&���{��n���R�-m�MY
 �XX�6_w��Giܔ�6Ȏ���p⻪kzc�o��Q��M�93'+��w����G�.�t�=��y�&g��x��w����,��n~�T��d��N%�P.�:��Ru��]�`�4��tc��˗+-(�[[�	4�(���-&����k�6�����G�P�E���B��<H���J�U�������I�ǵ}���=C�{K8;#\�ח��Yc�e���ՠ�syT��C�O��Li읗33�_b1A`�':��wiLUY_#�/��Z�W�fŘ�}�y��Ow=W���V�ebdI�LҠG@��j�e�m����
hN�\N��TH=���?p򊦶��LP��G�jz�9��7��v\GN��{�*< �>�`wL�j��5����d����Ȝ򠌃��
��}*p-��SϢ&+�����>Rc3�DԊ���_B���0/µ������x��>���Ja^��� w�:]�P�W_6�hʎ�`�p8���w��;33O@+-�{����5u��2�i��c�����c��9{o�wP�M��1���ጣ�"�=y�2G�҆}��_�]B5��'��y�O��ZL|�OEz��<�%�fS�r�������goݯ��ZA����3�M��aț�>e��h
��U"��ě�"i���h��b&���u��+\�Z6b�кS)p �� \K�ZԄq�u:�䨔�Fw��v\|t@R�'�9x�_`�_y�����~��2�=���;)�A�	�Lj/c^YV��D�e
Ne�B�
#�{���N�A��0����Rᇮ�~��lS?��
�U�Z������=r�J�r�+����w���:��gu�<)���gW��f&��pM�I���P�9f�֓C��x]i^hU��bF�f:�����Mj��j����˺Fs�'����i�G�d����1Ƕ�d���5�/"�)�d�UZk�@�	��Am#WK��u�)��x%ծ�%[W(o$��C�Dd�&};��8��#J�ݢ}ۂix�]�d*�ǥ�Z��j
a&0�<s��u���m�9�g�����A4śg`x s�c�.�w{6�Ut��#D�zo�R�7(�C2��m����_��{���xeLΙ���G��]�D1�|�X�M�6���:�c���/>�$��T��j���(
�u;��R?�j�`S�iA��WV��@Ś�Y�F̂�Sm�%�V����,Hj^�,#�A���cV�_Mi�6�0�Yn���R�[�Wm�9��ZE�@��[ݚ�Aʚ3:�Ȼ��&�l:CC]���e"��.�B@�i.��\�Y�Y�f�i0�[-%u&ƫ��X.�1c[���5�Yp8�X5��X\�]Wk5�nH�m-c��^&���Wl��cbZ���hZ�2͝�7���}m2mät�4�n���[e�i�٥��b�s�h��`)B�Q�-���{����q�Ԑ��{���'�D��.����}D��W�u��5�N{�T��ۢ�$R{^�./w�B�(�*=u�u����J�K����(�a'7&�M{��I��vJ�*���3�����H�����N4����t*�:3H� F���tӮ^���S��]dȹ��k�,��^��>ݮ����G�k3d=j:�)De)5���w��T��彳��J��1��]b�ܚS��ڞ��'!�(�^뚿�T��h�:U�݉�;i�3RW����! ��Km[L�_� MI:d
Y!a*��
�+��?�z��Єer��߮�a0"Q�啕����q�C.0������fnjcbh�
�NfJ��������!�@�w�v�>��q�/�Ue��h���+]���c������ͫ�益q8��|�xLM����x2Ɯ� +^��Ͳ�76���w��^��kO��JX��qA�1
�&��Yv̄Y��I�j@��ki�X[J��,�,�ie�U6Ŵ�6O،����F�����I6*�R���U����E�~���/�~�+8�o|UL� FM���E��fD^ݮk
ՎZ͕�޽�'*�M���lWĻl�����1Әo�9~��eu��o�a{}�Enͩ�_o^Yř����w���f�m�����6�+u��V����T�&T/�K8�7%Q�N��LĐ%z��,}�X�:�a���f~`�C�-����|T�	��h����k;�5e<�`=�(D�����6^s��r�@��D������_���3�{�+	8<�L�#��)j����C��ו�^�h�t:��.�����k���6��Q}���BH�^N(Bz��,�B�ܪ�*U^m�2^���Ĉ�垛�nǫ�~���仼�гܫ��*β-�6{�~��/@ཞ�:�|�t��Kr|�d�B����sz���J��ۀ�*
^-CQܹ��.���#s�|lZ+��x	�=5�`[��}�q0�eA����<j�M����x�t<�{Y����ڍ���/2,E����5ۥR&��֗Sm�z�b���3v.�\�CH7[X�]����H��|�mL��I��2�(fX�u=ޘ�=�'C�s(̓��sڷ.�R&5 ʖ���Y�j�NzzJ�1���y&r��)=�z��O[h_�7;���!���4) ���.��kO�Z�t�+a������k`�-3�"j;s�EZ<�}65�:��MOqz<��e6sH��L��[�j��ma�F8��*:�}h�9�<�^��[�;�ꏷ;�Y�t�6��3>��&��\
���U���ܧ�A�G<��fiu\�[��H�c��-�k� f%�zVs<n����ݟ���ΰc:�9���u8ˋe�ݽ(�^5��7���
�����X+#\kt��彍d2�@���i�����A}�#�d�rX;5~���W[2������7D�فϦs�"���*�'W�*(}e��w�}f���i�;����{�/a]�ޔ�+yH�%����s��"pVm>�ZrL��_�ݯ[]�v'�������U��SS��s�q���`�6
�]�V����c�7�������v����4k#��"�ymS�<G����0����� ��&;-�H���\ ��#��u�C0LgS\V3Y�b�,ф�˙�ᆕ�q<��3Y��ռ]�Eڇ��n}m��늮��>���hGl��=*������aZ�S׾7ً�\/�x�V=.�^n9�k�mEAћ�b^�X1�J�}��=~�{q�8��z9A��>v��5+wV۞QQ`b�7���g�������VI���M;����oV�/���%�g�t�$�&�EBO�{���3�vW��w�Ҳ�������9��������g��{���vZ���T��Q�2w����pB;�,$h�U�9K
0p
$4�ݒ����#ol��di3���ō)+.2�k&�G�^9��1S�0 �i�{�=�t(d��w	��u��ޮ�fk�>N��P~�ݮcz�*�w����]�[�*�������]��K0��3
�9�"R��.�X&�G�"x����|'>��Ž���6Ӂ��6�&��'�o;L��4֞#Sن�w�$	�h���#Kʣ�n{=^u�"�|��(�r���	rޓҗzz�q�G��*.�*Ţ[�p�)g�ц��WYVg�Y��JA��9[��`L]u�%�4lX׵�f$�ųL�s��][;��G���W^F\ߍ[�w�&Ɇ+/!�sEiF���r���e��Y��}۴����EQ���s>~����������O={M�w$�#$�g,�%voC�Ӝs�tA
-K�Ɋ|�Nb�p�[����/��om�O�"v�����b~�(�'ԏ�ˤ=��sʧl�,S�a(�������緉���/��M۫�C��bz���*�����No�d���sQ���T����ܫ!��x���b��A�Y�h]h�wո��򀧸a���;���67�����������z&sW���,�y�����i{L�g=Hm���-w}�'׮5�*����ft(?}@��Jb������A�k���_�~���%
 �;3����Y��¡��-o�}�z��������z���b��R��K຦
}��q5�s0 �/I���9Y���ɪ�3Qs����ٙ�S5��Jp&��L�M��4�Hl��ͼ��[¤���6��
ٹq�w)��eZ�"+U�3y���4]n8u�1q;��w��ҜҶ�(�;��nvɓ��!�����L+2��м-��X��v&�������6�ehWZE�+ޛ�q�.6\ǂÞr�E�U���ƍ����7
�m�oN����d� �6���u�;0(��Ku7�XS�ʉFU!�%n��
���7[�6I���W7l=���"����uo���M�;+��o:�v���*���4���}�R���5oo�v�s��X.4:;$=��	�Vt[��Y%�u|z���X[W�=���r���o�>��C�;C�:V�>	ڻJ`��ns\z��,�;�v���/7��l} A�:�Q�koh�o5�.<h1f�> ���׎�����T��<or6����]˼ꕰ��.�v�ul��1��V�VSe�o����gf�T�/:s�Ayg����y��Wu��w����DV���G�E �9��h;�]�J��$D�,̩���	u�e�s�v�]tB�,C/v��޼�f�I��f�_�f���j�v��ݦ�WQWWY�����=� e������"U�gU��ٻ#2v�g���+��_+��v3r�ý=t��v��g.w>}nU�yՋ^Q3����͡�u2��7�QY�@��fg���Y�9�;R�i�t��@�xC��f�����P�k(-9-V�z�L�����9Vl�
Xw���o����8WrvO;�a��5ۀ_*4�koL4;�d*˳\���Z�1� ,�&��cB:��q�g̈́t�A�K �u%���`�3	�)
X�.��p� �fq���	���S%u�Ff��W�h�-���h���H���35iU��E��sV,td�E�4յ�ՙě-����d+�����chf�#��Tp����6V�Ж�!�����풌s���ڗb��Y�B��1���2ֽ[-���%î���7ie2e��PU֕�l���x!��L�hb^қ 1*[׭��LAL�h�Yt.�Y�C.�e]]6�3�m
�M��i2݆&`-\=Gbr����ņ�І52��kJ�1���]KT�5�hj6���*^��\��U65�jG�³bғKR�Wu�������څ.62޶.��\�� �m�g9ճD�,�l�Ӛ`��q�nF�]li,��6����sv�BbR�F��]^m��jЗ]��j��p:���v�D�TF�hb+J0�b�:6و��t�m��Rmir�ͫp���M��լ\]C�f��襤�b[��3�[ٕ��󫊎���Ghͱ����6s��u2[���"um�iY�v�bԛv�lGL�Ś/XA�hݚ���s{K3���k6%�.&9I�.MK��&BR�ö]��4s�V�e�Ԯ�]f��n-f۞-Yh�A*�V��ޭ�v�V�麗�Z�[�um�[��ݶ��BZ����\E��)-W,׫��cJR�Y��m�s&��ZZ��#�<�F���kkd�g4&����Kc31�f�p�k6��6��f��VнKoa��hͮI`��k]���iqq-hJ�pYu�3�q�q4��5�v���[Z��[2�mjj*h�f �˂�)Yc@mn\Wuq4��h'7W�l@	lFl��F�tB'9SKֳ;9�nݞ�.��]Ʋ�vF��d�Yf�[R�a��&��5��
Bhd���5ͻ�ļ�h�m�ZG�5��{Z�1+�V�m�i��	�X)4�hR`ȕ�ٺ�(�	2`��*fY�BjR͘%�v�]`�-��J�@5	�#eH���i��m�݉F�L�m����;�S��8$���<NwS�����+�7Z.�chA6m�%ض��6k��2ᴵ��\:����e��٥�tfHa�K.�n*��9e
�6[���:��<�BvЄrPғge�#�r�)�VXP�]Qڵ�m�Y�b4�%M�)-�2�5B(�!��qK�h�ջu���t��ff4%���`�u�7�jM����m�teP�[{K�Fٕ]���a��[y��5\J-�4]�����V`,��)B�44^��5�ٙj[eA5p�a��`v��%�͓&5�K�q50�o��#��z��QaHخ�7�Y��]��<���3޼�@��ں�B�Y�w���s�=_V.'ӏp�m{��h�w�Ь�!��O~�ĳqwԕ-�))h\u�rQ�h��������i@�M��_u�j'�v"w����ۈb���&�j��r�����]ei0e���â�g��E�<Ll��m�VA�Q�7ǭ��F�*0��r�h-`R���Y�t�~�9e��2�Q�{7	�B��V1�F��x��H���T+6�ûyZ*U�����=��FA�Qe���m�в�]lu�C����.p�z�U�U3������Nթ���Q��jȖ��y�߰��Lnt3�/�3^����t��m��p�d��`ЄSM���M��r�mo������x��u��BYU�x�(Ӽ�=*׫>��h*���§�="&)|�y���D���bb�]S;�ۻ��{z�,��j�G����XGL����u��P�:�`�uXn���κn+cf�a��"�u�@��hڗS�嘌����W��j�TH @�Nd㚻Y/���4�ף�bf���;�|��	��W�[�Zڌr]V}��ϼ�GK�<�_�L��j���'xK>~�T#v���f���sU���U��]n����ޜ5VK
��c�]�ֵ�j�]��n:�B��4�W`�&n��5��w��p��Վ{$�w���u=��=m�0[4�����x^���G���S択��s���Bc����#�|���@�+f]ѓ��\��k�3~����1*��u�^_֑���mL��w��X�E�&a����� �a
5ɤ�v��n��8��>�>.}��=>�џ2�
w��h�%!�_r�fd��ɨ5@����)����5�?d����b0P�U�a$S��!��[�D�]��c9߾��B|�z0�Խq��~�6�EK��:qS7��%��uj.63%8s��)��T@$cR�0���P=xv��U�a�B���6�h�����(�i��eo]e�[f)��2�-���y4�2��Z��9���Cx�r|b/���SQc��2(��;^�~��XȌm-���W���������H�dy��u	��}͵E/k��<n���(I[P	d�/������>�toy��|};}G����@�ϣ;mD�x�f��|'7���Koߑ\�V���n��x���5i��_�|ݣ�G�p��R��,�(麻�?aAx�U�|O�������>«;�����:��\lQO�X�t�.9P����I��Q�%�1^�UM]�=v��7��k���)�fl����0���߳��Vi͵������'��h��Y1����������%5���S��p��/sՆ�|}�t�D�UC &�Rq�u�:���(<�|J����6�����=���,��7�8��p`��&��7���+�Ю=��:�n;��(g�m���n{r%���ޘ��}>�Vhu�8�qL)���
#ہГ�U�_��Qo�W/�
���χs�)gzθmsneU��-�@@�`ӓ!�-Y�vk�l�a�Aɻe�Yl�+fnHb�DS{�&�����-�xg�������;�g���Y�e�ݔ�f�u9���:g�3�
F2g7_j���������ﱟ9e+��%g�yr_+��LA#�O�[�`&�ί'�F�x�P=�[(����#�S%f#yf�VJ�
��yB<vo����r���fL�[R.�1Z[c�^��o�b<�>x��u�(2��-]�&�޲-f���_�f��6��K������j����>�	������V�ae��8݀aq{~3cUg{z���w����9�4<<$췽>�[��:-8U���n��&q����ؽ��U��ل������+�,!��� ��^傧�o.�^�}�Fn�e�z�ڔ)Y�޿�%+�7��͜An�63�e
�Q=������6��Vz��x�f7�y�J��`� ���κ�����B}��lh7v�MV�U)��=��Ꚍ��;:������Y����qRr�P`k��췧�"��,�(Lm�
c�cӦw�� �v��F:�v�a��KA­��mXJ)B���k�U+ Z��M6�m���������M���s�AI�d/Qǯ�qB�w��������@��]�~Ƣ�ߜޝ)k��G��h��X�vU	C'�x�4HI8(�Sm�b����.κ[��nc�g+Ϧ��7��06q1���T;~��7�X�}�����8�{��_��ﰸ�?{�W-1靝"8�GzPZ�AO�)����,-�9�ם�S39z���@m[��n��3�.���\�sE���U��`�i˚�g�<�U����ѳ��µC�݋���E�t'� ���L�[W4yif: ���d Y�����qף�
�^㳯�툸�C.<�G��=�c�x��}�g�j��%���.�5��N���I#���"�JL�����m�*�^1f	G��2!�:z��Q�vUs�S�����r;\��W���!�%������չL���}N�����f�l�Y�y����ȕe5.�;�GC�vˠ󉙣�n�Y�@ͫe��3	i�������Q\�R�Vr��Y��{��!����#r�k��!s�R4Ԑ.Y�%��S�Jh�F4D��Ƶ�Y�"89�na6z5NŌ�Pf�m���aKv�M��qG36�u�G,-��6�(W��Yk��k�jP�͸�-�Ұ0@6�7\qy-`���@-a]Ś��*�,m�$�E%�sv&�F����qH���ʦ�k���6����]M��m�D��\�7m.�uRF�!-CB��>�����Y�mf�l�U����D�b�k��un���5���m� [�Yh�-M; 7h��u8!B�Rt��<a�b����|��%�,�|MϝP[�Ɠ*�o������ W��p�5\*���7h��!�e0n$p2f?wa�ݵ���޳��v6R���#�1�{�uș���8`��4��P�0�%��}��Q�N��z��N;]�)-���>��50T	�]��e	u�ij�n&ޚ���/�M�"�����-�0`H�'B��@>���]�^�1�,�󩩖|����I��̯GWV��K����#`Y��g� �"�4A �>G�ںr����b�/_vb��`
�U6�v��꟬�ټ�����PĮ�U���s?k�]G�:��J���in{��grL�U^x��B�BY��9�.�Z��g#��jp�o{���n<���Զ��%���@[�m�t�-Pۮ��{��y&^��b�'$z��F�h���U���^b��EO����R�(#��������i��&�P��P�]{���B�[�5�i3Y�ݿ3 ^�eB*������ViO�����gH�8v�����_z�z}Fi(���q��jF��[ρ8����P�<�_U��bh�x���T�j �%�dYnξ{W����
��}��8v�c7`|�׎B�f��E�}�\�[
�a�N�ɍ��bEұ�-�Nk�I|N;yB�^��P1�_pfb�b,�E��yl&�����~7�^3�-���b0�d�:�"z�g���%�8���<wp��_����U�Q��J�ܽ�]�����5�@@=.��n���q�p�G� ��������5�Y��^�N�ۮf;;g=�}}��gW[��T" ��P�ooȻ�x���s�c�7#��Ԡ<
���ntxw��o��Ģ})A�4xڵW0�s�����Nln�i�dn4�7<�˵�k�6&7i�a[�i��N�!6��Q�3�����6t�ߍ稙����'���r�W�4���M� �&L��TK�$��დ�I�ܝ�Φ��X2U|��B���KxX��3lvt;76R�/6km��Q�Q�.�Y����퉁5+�Oe��W���1�Ob9ݷ�k��$V�`�{=�/朿�*2�g#0��7�q��^�~���C�ޗ_;ѽ����$�	����4�1-S]�kG�=�t,���ueE�WϾ-ۥs/��r��ǴN��]
Xe�;��\^��{�}�ܷ���0�#O���,6��2�PQl���G�'�=�:O�o)��:Z�]�ő vT��XNk�J{j���Gٰ�ڳj��]|zi��Ň{@�VVѻ	�o�mҹlgY���j�N��u���ۗL�7�s�zճ�t�ͼ5�-f�RI��j�ﵚ�7;;T"p믗e�{����r�g�n%~WW��d �d �s333�Ȯj�-��
F�K��oT|3s����'�{]>>T��F$t��ິ`�2R��r�`um���W^��ٟn-w];�G���qI��-�6�)6 #m+�`����gR�1X~1���k����zj+{޽�^Lߏ��R�ںc~$�$��5GRng�ī�3�I�F�[�G�*����0�����"�V�#�)Y��cg6�f��knin�8ְظ­A��A�k/�\��V6{�٪}��͙h<�:��u���[�����z缛��q9]�7��$`�w��k<
\To�=���4�>��(�@J]糏���PJ�U��?q�8/b�}��Oj�Ӝd�ɛ�cԓ�
������W΄K<�S}�O�����389t����H&�#+�Os��ɹ3������$P\���)��f��4^Ϯ{l�':����7�!��*|��~��Lƕ��sgЇ�mr!�UF��Q���8T������6j��q����7HW�$*��5Z�8Z�y��LD�+';�����^<A�Qx}��.K��.��-u��˜�gUYH��=�ֲ�l8NV�u��#;-�qSFa$mgp�w�����Y�dWWG= 9���G�)�J���1���V]k�Ý�����p�X���
B���ߏ��̎�3��z,爓+e���=��H�;˙�����u�Y=f2��@���������{��,1S*�}�G�w'��3s E�X��J%.�5h�YI�م2׵75iq��7�QЁ���.���Bu�TV�Н��޹����:b�Jsf��&����0�\���Wq5㫗�n��O�|Q��R����ߞ*�s1Z8���|f����-�"���V�G�������Y�$ʑ��a���4 ��{��+�����zd��g#z�8=gG�9�y�έj <�ԫ�	��W�L \�x��a��@-�we�_ag�3�g��e���@/���7CӔ=��Bp��M���}��e��aTo~��%��hM���+J8�; s\�X�������򪀳x��%X��{�Xn�t=��/gܳ�xm��Ү=3ȜC�d{|%us��֟%.7һR�GLd72�0���X���x�g�w]E�Ԍ�$���u�J�Z3X�z��ei[�T�h_Ūg��4��	^���HAp��������&���9�Q�m��(��$�WZ�G��C����뎃��:������Z镓���q�뛝�`�<�VC>�[K(�
�s���&��SZ̒�tЃ���5�VlQ4fk�X�0�٠���FAwR m-(-/k���LSK�n2��m�&�e��K�cZR���n�%�+
�h��˵�gRd���v��]�4�J���\�\��n�#1�qcP�i(�$nҦ����b�b��A�d��H���h��1u̺]7f�J�A%�nff�#��VJ����޻���G�K4лF^%�M ���Z�F�(���	D�4.�S7um1��5��2�[��&����`O��8�3~��Y~�UkhȮ#�,̿s��o�[­_�i�Dx���z��E��Lxd�9~�gX��E� # P��\��f�Ό�{���0���s)�(E���ޭ3+��.�E)C;�ƻ�"0m�a��3��=� Ny|it ��o�:��iWZ��J[E�
�@�}��{�WxG��/�O٪�]?ܠ7_K�Jb{�z�GUW\ma�dj���~z
F"4��>E�;6��> 7pd�l�eU�D#	��f���l{�m8"�? I%����_Y�?�/^}q�6'���>�-?�q�v�j��U"ӹ���3���Ӹצ����� �iPnfb��H}�v��ۥ����y*���a�M�UT���9ݟC!�7�;S�N���q�Y��
���Q�T��&��{/<����Ok8�n��\kd�暎��7m�j�]���5�����R٣�ݦ�u�C`�,.�J�D\ ���mx�˙_3�O�3k���͈I/s;�5��D�G�������s��G�|[�8~�S�?�g�9��l�4��3�ί(����R��@�0�Z��[^�me�;x�x]���Fw�v���n�pʣz��&Μ�id��B���(u���Ch��T�_�m]S�z��Wb�+/bC��M�*D�x�hѺRh�������j�@>���5�g�.y��uQ�J|}q+�5X�kyw���:�}��j+�`�jE��Q~��ɴ�E��b�<���$>옡�V��R����a��/�>�T��Ծ�y��88����W���3�':Q0�Z���]��*"�X�)1����N>6�wL�}��}����������CB;j��_B�=�Re^8uW�fj�J>�d�ݚm����۱��ۆ��.�4k�n�	�_|�QIX� 3�^�~�yG2ۦ�����ҵߧC ���0쟸{���{�ߍX:����ֹ�as��a@7�΀�ϓ$p3�o�I���O������QK1�Y���E�&@���[]n#L�m(g���-�%Ҩ�j�JM��HN,���
t��,�ޯ*�ݫ$��tzjusه��Oi����ǘf���3��>!侧� "�ݏ_2M=��r��.�+ҫw�p�K�m��H8~Ǔ����fFP�~༮��G'�Q���MA����J�vg�N6�9��YS��c�B�Ԯo���H[N��4�O��C2��N�Vw0
�0M���pӏ�y���	��g8>}	���CŽ��N������,�ݷ1}�+v|M��ZB���h���O&C��f�h]tWV��eI�:(/������iktm=��) kFI@!����Q�]r&�gfWF��S��wC���qU�"��3]oJ����"]if���2fMj�ۭdJ���ÍX�ۡw�!+�/��	w�1a���N�?w]���sꗇlnٹ[�x������Զ�t\܋E�ڊ�K��+%ҡ��Ζgfe
5���m��F�|�๲���kx_��1mn�G��f�s!.�r��p�<��<��"�E�9�P�rŷBT��5(mm����*ڷ��<�P��J[�\x��ݯ)={`����B��M�����$*+�α���A���g]��;�x:wX'Mz�V�����M�ҫ�N���{�Чa�J��b�r�So�)Λh�Z�j]̽����	kC�hV�d��;�x�,�[Yy"M�l��|!� �o�,�t�1��ۼ�Y�yF�e�oN1���]o[8�N)J�2K�=XTޡ.����&��s��M�U,�������c\:�E��y8\�,�IVe�T�u�G_V�EvC��]���V.۬"nfe�����IoM�rh;�-:�6����]�̜� .90L�TcG�l�7��ͨH�%�Fg�F"�F��:~������C0i=��Q�˳�;�c
��Y\VX��@����z�\��W}�vn�<[��-��iC�Z{Qb�=0��B����z�+&���E������}��?���TkT�k۫�hйݔ�w"�c��|P§q�p�<*��w9�)ߌݳ#��CG�n��7ޟ�=0_c�|3��Ώ=o��;�p]xϷ�&a77(��r�����1�f�I6ww7V��؟tyJJ*M�A"���T��ָ^���Ɋ�K�Q�Tϵ�LN�q��F�;L��O�����޺���T�r���u��C{���h��p�]]|�zR�>�W������\�U�G����^��}�������A6��y�U�<���m5��[W[&�n��Weq�����ppk,��7h�v�HH�d����������'Zb��j>�~�R
+���d M�C���gp���n��Y�9dEW+�f[��^��\�J"��j�PZ:-k�{tk�Yh�	-�!8	�ꇪߦl����)���s�n�r_�dv�:�!��*��؁�+4��������]:Z#�*�)��5����Uc�3�>�'�m��n��@Pe)s����r;*M=�uŷ�ǒ޾��]��e��mT���M��s�<����*�^��y�G�/�W��>�0�K��>d@�\�M<s���J�]n]���J�SZ7\�Q��Y1P/��+1f�fh�;�*u!�d�9�	��k}f����a`��m_nN쬅i�&N44[�@~���9����KE�s�f�����6�Q Ij�y���?�׿ui9W�;-�������ɞ���ҭ��m_l�������o�ۻy���g;p�S�PzQ���GC�3���y˜����t*�8�*�Shc�cEz�N�x6ƸMk{�9�ν��OC�SC�Ґ"�ػk[I]�X�Mr�]l��[mi�u���!,x0,\!��Dªc�>����N��>=m�5Z�r�p����R������{儗�k/�Sy3��K���W�"w	����Ƽ�G�~Z>���3�4�l6�I���Ɔ(���~�W�t��/�sQ��Ҥ0��Mn��HI�î�?l:�n�O���$=�����m���;;gO����ȝ���N����`$Z0�l�oc�j�a5�nT!�Ɏ�d��b�wf�B(�]Ta��tDy��>y�b-�.l�����Q���k���D�����3�5
��\~!��dB�6�WJ���TN��P��.7נ�®���� |��4�
﹗�fJ���d��}���{`��5@�ױ���BpЬ�m3����E�w0�}ٌ��ܱ� XFC-�n9�����ȏQ�=��{�c�@��ک��Ղ4��</4�{�TV/��J&<ls��^�S��;=Y0���n��=�~u>Y���#��$����L$��"��Yp.�&<����vR�~DJ'D�0L �F݇p�)�d}k7o;[��RH��3�Ϋ�#cB����1]��[xם��i��	��,!M��-D�ͰYu�D�d{&���6.]LB�q,�+�����J��YbZM�U[�F�i1ZH.`��I�m3�U�k]tK��V�z�]k#����6��!n�,�	��ve;1cu3��lt5��]
�m���hU�2؍�T���A:�����ؘ %e����+[{cn u��j�j���n�-��7X �l�1�!b@��,תJ$Q�����(I�r�25v6d�;��6��lw�y����Ey�4)�{��Z����׺��Z<���o���'�2�K�W�_�}���.�����rp�][�uB
�R�\�������q�<���d���۝��� Bb��s��8s9N�uI��~!�@�P�s���~��GI]�r�e|��c "�F(�� ���rq9��7��cXsY�.�g�f�N���y�c�yb<1g��y|��������Ӑ¥wfx�*�>SA���}��vì+��42�3�W9��;�Ǣ�i��Az8\w}&�����9� Y��7�=g�z���^�Ue�U�=*{P�;�Y��S���@��{ޫ�i��>�	"�@Ap�w�vJ�{r��=W��1�5�W4�^�F���KW�~�T�kN,p��8{��0�{�G��tn���G�^�
��u��a>�5��y�M<�ɵ
�H�L�{J6�+sk�r͈�Kٷip� �0��F���Z�cp�RYS ;�{�7�Tziִ]g�͘�q�7hyﰞ񸞽a�h�����LJ������2
�z�S�N�x�v7��>���ut��ư�]�p�DZ�+ �5�,�zy��ٿTX�ы׎�=��>�#ꑘ�����բ���؅�4h��Ϙ�%D,)j����؎	��ҔM�o�ά��`��� Йu��#+\���%�]1g+W\���_k�������_���v]�?�'=��~�Ao�c_ǽx%�QH �pwq�����>�T���>�p�'�0֊z�_���op�N��=`K�97w/;%N���ƕ.�5�+��D�^+ﳁ�g;�ߠ¢�D���� �a��|@��Fh�{X��ǍWR�����~���"F�Uֱ�/z�p�H��{w�8�-��p�\y��0�f����cX�k��`J�LB&�t(�o��+j���J��/��n.6z:�ء�lL��įG��I@���\���\.�!�Օ
��E"��{M;�G��$���>Bp�J��`#��Yi����)��ls��v�s\����-��ŃY�i&��WK}�k��N��]��XJ{�i�^W��w�|R�gz�|r������J�g����>�
�v<Uݪ���y2x��ޜ7�Ѐ�(3"S�����5���'�2{u��s�>�Z�҇����5�./+|�E����/6��*�!	E/��ZI�k��+����=�9xw��~jd���� ���"�%3w���>�ۮ3�����h;�)[�F[Qf������Lk�u~�Q�9	U���؅�aǜu�ʆ��kn۫���e��th���hlr�v�U^�}�N�ᇃ��-;i�Dso���b��^:*Ǒ�����ˡX&ZU�V�$�J��E�7cI�`z{�rZ�
�vi��5h���Ė�Z�T:����w����"�����>^��^����|I��W��p}=��M���' @.oJ�7%�St���ɍ�= �OR�'T��|���/�x�鳷�$k�qX_,���uW�٫�p
�A�����r�\3$��?o�
�s�-w�qi���i��Tx��]�Ɣ�9��S[����r�ݶI�ct֌s�X� Ai�Sg�9�k�D�,�t�O����x�f��vx(<V�g:=G=�B�֟��}:�η�AF9�x�	�X��ڍ�<:L��p(��Xi�7&RE��`����n��^9������}����t5�{�t�a�"7�{�%��}^r�kXFi���&��^�A8��>�.����5_�+���L�]_��&Is����/E<H�xd.v�Oz�&4\�5�  zP}�6�����(WL�}��M�U�&[���Nn5Hux^�^�5)\r�z�lr1y���P����U�Ƈ��#�@�����@ޟc�c�f:��&ѯ��G�U�: nG/�� +��b�8��v�����ۜ];u�Ӏj���n��Ԫ����G*������r�U��~��!��~uר��x#L�k�%��W!%5���ig;�Lō{6'a�"-^t(��1{��U�U�2j°��zt���MT��S#�c�}٘������s{�^v��;4׷��.��F��ZX����k��i�Yv��K�3]�fc5���`� �#N��8"��qJ1�[�>I���`�_�ݙ��y��z���r3��T�����䁛�s��%�,�Rl��KaOv�'�ܵ{MNV�>a�6�L0Rno����P7Jz�>wo�.�CB�]2���85�αU�9���9��"5IO8w�x������5�s�z��o����h�ۿ<]3ryu�ݒ7!#9&k@Ų�?J��;���tc�9N*t^8�>q˖�k�������6sV�>����׽��߽q���F��7�U��s��m*h����}��}\�e�Pk<�1[�֮�~G�s[��o��f����?�N��������=/����K�i�o껵�;�\�;�,h�s�d��TT���L���	t���v6�l��Q�����^��cC�U%C�z�D��]y.*	��ʮ�ѹAX��덹oS�t虂$[3�~�"Rw~>��v�D��dŕ�qF���g�N�)ts3!�V�{Ӹ� Rw�3�c1���3��ɻ�9�+��j�:�E8��Ee�0lrXi�n�0Y�gV�65�=����ٍx��q31�q���P ��d��E��&c�)���4mqh�7��r���i����n�@ʃ�k��-4]��G\s�K�G8�����v�-Ŧ��1�]�k
�l��R�#�L�2L���n�nnc��iJK�u]��͎n�u���J�t��W�i�����pʷj��?��'���RK���l'���"�nЋuU�d��;��H�K��XD7,�F|T�{��៻qA��{Fm�h��E�^��b��e-W�La����=��,����3��D��v;�N�	n�:y�3w����㤔���Ӕ[q�LN�^�sc�O[͉��w0#�"$+���yP�$Q���^4_Ug�+�0'��=��'9kr8q/���Y,�yH2�5-����r���uݲ���j��l��ǝ�8�{�<����Z�]�"��J]�V*��}0�N���WX�N�y�,���GBh��
i��P�i6�+�Iǌ���3���9��WmQ��}JMS�"�&ΐ�,�zc�!m��7�3�N:�U2��}39����u�>8 �d>��zǰX$��˄�2���'�͇��M̎�Wș�uz�;s��Jh�:]>y�a��P#��<��ᑢ`a>����~���1^I��#Z�y��r�y���ڜ�Eh����v��k�I���7c=�б�t`��y�m3Z�L�]�3-3�U%c63�:\��* �z���w�ٛ�]�o��(��p \}�s�\TԄ7$o�$P��;�ꔢUM�3�[{��&�P��b��G+E8��UYy��gA��۟�4�7`c�I�b����`ڙC�����˽�"��e��g����}XE{ޏ�i�8z�H3pc8�ٹX��o	>�eJ6~	t�kS�Ɂڨtf{C���3�'U��cy^먱q�p�m�,2fỈ�"�ۋI��E���2SxNb��2EWJ�+�x��{.���׽��y����F�o�9�uE��ֱ�7Z��S�G}��m������޵u�G��M�s=��~퀅T+J�6��)�7�1_;�%�=,����!V����M{|�&}�p��|3�j{0����z)R&߅���y�_:=��+�N�My��\�{AUb��+"q?Pї#_u���V<Z�V�L�u2��Qs�;��m��a�x�Z`�8���lsP賦}R~���4R�`>O�/����osˆ����Y⥂vsu��Ԥ*뀰��C69�k����.���͊DFP7Tt���_�8a�㓾�}c���
�4�u}��w�i?���u�Ӿ��`��/�TE��A�>�%��}��v�����`���:�"��a��u~'^eaQ{�k8߷�b��]y�EF���}�UGT^�"��~*n��+�G��G�0�݆���x}�5q���Ύ�����5L
�L(g���k�
�eg���Bfƒ��H�ёFz�(��ok��[����R�Zz�g�P҇�X���⾘U�뫻�yn���Z�sC�j�h�t�A��u��>w����ߌ��I��I}\�븛���Ұ��q�m!�5����M���/���=u����3��?]r�c	�T�w�Ϟ��𹒄mwa���Y_a����Ck=��M����.�0={�XAd�2�W���8>/._����;�⨵����q��@݇Ύ�m����m�C�V�O���9z��p��T��o�bI�>T�خ�|\
�k
>W����O�N�ci�|�����ILV�ԻZ�1�2/maUv�[����Tm�ۂ�K")��g0}��#�������z7��$)��f�����aD�Ӟ���`Mn��d��z2�2Ȟ����.�u��}�:�bȹ���N>����ݔ�%��l�ۺY?/IyQ˱T�ֽ9@釳x���^ij�+r�w6G6ϡ1�O�ױ/q�y�dofa��wB��p^Փw~h�h����V����S �%5���Q���3���v��)�5�X?���s�8��k��nI��lzGf�U�<7�7W�`�F2}$=��Ҿ���H��	U鉐�ة�z��L���r����SS�������⦧����x�IC�����{K<�.�I��S3yu�R��[���*k������O�O1~~���Q;�U)qa�|zE�m�WJ���L8��AXj;k�U�;2p�`����4Ѭ3��Y��`GM��2�w�t��Cc�q��*�g%t��{�s1䂘����� �	4XI�w��� �j�+��1�٢��	��3*��-г��|H�T�(�X�Jr��3+=�qU��y��V�=I�^��=7�����EY,ї��g�߾�.U�����eW��[�R:�^ל8�Xe��.ˮ(�R2�8����0RA&���Ħe�i��*=	I���H����,�7������N)*6eC'-���$E����nr�$�����0C��a|������͈�ߪ����B������с �ok�봮yШg������N�=P��7��H����47V�^�_NF$���40�V���A:��c�t�'jVϐD�{��
ifN�f@��(AJ$�<�<Y��hO��>����8����'޾�k��s�h{��ݪU�>��h]�Nv�e��:�Ysl���D���t*������z�s�B��{=W'�+3gYwqO�n�)��u<�&
48�w��z�`��Iq.�����&��.�=1X�},������քGe�( }�\M�B&����ӛ]b��FZ�D�@����j`�	�lӻ�).�5��[����sQ�lu{<�'2�d.:�� �h�:����$g.�Q�"Ÿv©���@D�Wu�5\����,��g^�-C/+V��}��ޮ��9.��gA�M�WzX��M��n]��ŴFF��ė�}H !\����2�R����e7�v�L̾{�]lS��:�P���Е����`ү7X˙f[zUe�mlu;ow:�w۝�d�[n�G�'!c���Nȯ9�bE�Od�Rb�ǡl�yNP�5U�jǊљ�:�eA.c�ͼ���%�Ew�E���Kf���Y��9{��X�^�;)v��$��*����:�qɏ��7��aIJ�o�]��#���z�n�
���&]� ��m����+��V��վe]r��0�ͬ�V��4X.����/k�-��;�,YP��/)L"��� ��8��cL1*@�Nkά�6#�br���(�b��v\��W�j˙2�̽rq��pC��F�%��t0K���ݔ.�)�	5,K��]�p��Հ�c��oX�y�h.���r[dD�`������\�������U��/y�;B��W���3�]ު9���xLξY���؇_�#�R{�j�l�H��k���v[M&]��Y���~�j�P������W��)`��rB���sF͊:������wͬ�ϻ'���ˮ��]"�k��Ў�X����=suLn�;]Lb��K�.�X�j��M՚-Q������u�}�(`y���mfm'�|�l�p��+w�k{����sGj�7d.9R[��u[R�o{-��*�<�:v���[��.��阶�n`�W%)^S��[.u�8�QF�HS*���hL5��96鈍�B���qb�kΒ�@�l���f֩��k�Er���[�4����:5R]�7�kEv� Sj��V�r\�tf�3f�n:��ص�1tؚ�U���:���b,J�.��q,i�&s��@��R�[C�2[4Ե�5�	
�l+%i������ܙ���t�1���^���P��(�f��]�%-sH@1z��3;UXhwb�І�Θ�e�,ֵIFa.V�\�ulih��-��Վ��1F�h�Ҝ���cպТ\�[u�iY�ĩ�uU0�t]���m��F��k �dk��ٶ,�XcKA�K��Lƅu�͗F�y� �Ү��jٶ�f�l�4�m�k"х�	n�I`m��#�f��1��)]+��!�4�n��z5%��U��^�	x�`u��%-�myt��f6��,ї�eݢ[��Y]%�f64���&1Յ�a��AI��[b�PE��RlU�̥�X�\9�T�30k�\�������l�.l��n�c��	��5 K]���:[m��k[4��Gv�!��.a,�i�9�JL��jm+��%U�f��t����ĺ�����I�����+����ݘ�m�5�j�Z�t����ˢ��:��@ji�lKf�p�4�,ݍ.����b��XA�7M
k66���H[��`,�� �ݫc�b7P��L��K�ֆ:�[t�kH\[d؊]6�stK���Ie6��a3���W$Y��@un1�CEو%�,�m�R�;U�KHD�Ֆ�b�<�em��6�@6"m]3���΄t�df�2������֖�K`%�t�M�Y�vɯf�nn��Ў��3K\�+a�h�f����h=����6.���!y�����1�ƶ6��,�gB�5&6����n���U,��k.��-�aqh��p��3�U�%�"�������kd	���F�n�JBh�N-��R˷5�K�ג��+,JW�L:��7,f�-��V���Rd�3[�$��Z쩵�@Yx���@�x�鬶W5m�2�n˝�L�լa�C��a*d��Ɲ������s�|����v��4ň�sK� GX1�t՚5�֛:[��u�rK-�&ډ��]��u�a-\\S�hYn���)�qnXK�u.�%���[ub�)�Shbٮ���e�P��e�Gi���ݝ5�e�bkJ�d�uI]@��ͬ���f��UB�.�6��u�Mv�شb����pnst�E5�en�Q���h�
*� n
�!*�&v�e�m��.�ٸ5-%l�͸��s���j�^���qTY��6�Д!.Y@^�c��]єe3mj�K~��_����&ݭ�v�q�CG�3]򖼨�����3�ΪnϷ:��}����N�d����ϛ��.���`�RT:���N]���eS(>݆?W�ԉf�䝄Vx�]TL;O�zt��3`%�{�TM�]^�U>��0�"4F���]V @v"Y�ޡ3�[~���M<�qɹ����8ª�1�ɐ\��[�kk�B>���g7����%����ny�r]цT�r�1~�и��K�i���k�a�Ǐ� m�a�N�)]"Q��g�$���$nmVNN�`�n,P @A�Hc�]b�h4qB#_]���MQ:�ܨ���W�Tj�k���dVz*�_���3yɞ/o�) e�$��Y���O������X�2���ө��	�!w}�(�Wg�ރ�^����9��]�
��r'����H��"�r3��oVd�kew��-����l����]2�:ͥ�.s���f�K�)I�I,jZV�ԕW1�B�,���L��\����}��v*Me������kL<�1%���D%�jj��p�����́'I^
�! �g�`���[�ʩ8���U�@m��ClCH�^�g)�`
�1�s�X+am��Fk����أ&U�)&M%�]���x-���kQ]�����C/��.t=a���|)�f��◄���>�2��}������&��Ġ�>;r�����1S�.�~.��W�����&��=e@��W��B�� >K,���T��y�yrqȚ�#���m�f�I~�N9���7�F�`;��=미[����y��O�lw1,���d{��v	�5z��g�Xr|�u������e/��`�`�Q�ޅ�{�+7���w���0�v1�Ֆ�}}N����2Z��pt��\�׉$���s:0Zp��[f�_�M_@'ˤ���F��FhKjf~���擲�)[�ӯq
�Jt�����өR�g�9s�z�͊��gn�\�قp|��ӑ'��αC}�a�LG�s��bڟ8�t�"T[����jw�r]� �f�-u�e6�sn�c^mڦ-+",>
��h�+����9���C3gnY�u��߁�vW���.z�ޘ��z�ެ��"M�����.�}�*��uD�z��Θ����@�<~5���A!"�(jA�ٜ`�����پua����m��5^�S��j�7cR�%���̘��no��p/������6������yl^%]{a��A���)($�kǏ}dQ}R�6{�zc�yg��;�e��T��+�g�[���1�ҷ��t%��ƓE�88֎�S*�����#,���p���J��!�%v�ȷJ�S��1k����gj���Q%w��tc$xA�]�s�@�
�p�`�^�G����0��I�h�s�.��5+h���!}Vn��"�`x��s������Fϯ��K��$���]��Ϻ^:�d���R#�� �f� 
 ��ʩ ��f���,�ٞwݘ�a��"��=L����n&o���:�G�/S�Y���{��(�i��(���7�,mb�k�㔣A������%��SC){b�����ͭy�p+��d���&�HY^n4`��H1Q�ʂ�+
]w�����7\��A��|�Z������S����'Ô�d�)�m�f#,P��9o�ڗd���qfֶi�1`�nZ� � B��Γ^�ze=bgV} �\����(}�x5s��9M}o��Uzy�wM�1u�����6~��}�{iĎ��t��=���ޣ|�@��5�yK���EZ��Q�W���& �mq��4l|>�������\�=3ѽ�~Ed���g�P�6"���gf��L�Q%xx1/?u�ﰄV�V&x��G},���׹�w��q7~�\.��(){>o��aՃ��Σ�O��oO�~�"��3�|���ֈ�EB2#�������7�VNf�ֺ���#���0���͛O���8������a!�%�^����5�:�5ٳ�Q���?t;T�Cd�D��^SZ����g}�4"{8��g��$��x�E�L7�섲�(�8��Q��HU�d��H(�}|��(�HZmN��X}lǼC8P%����{K��qn6�CB��hƺ�K4	�SSK]cc�.̱i\�)��]�z��"�rN"���/΢��N(��ɘ^�AM	�.8�=~�mo/��|݉K=�
��G�&�c�r��QpDi��Q��e��k�@��f��ׁ�^�v�9ؾ�>o$���HU��b4�Gq΍rf�%��l���e��gڊEX���A�GF�9�UO�_Z\�T�9�le �(P��u)����T�r�Y[���Z��}�jZ�K9�(���u��*����D��d�?{������ظ��\����<�2�@( 
I@3�=n-��^��u/�5��}��U���aŤ��,`���L,���ߴ�����j`�ݴf�޲>��5^�{������ӗzb@H���ݾ8І�!8��+���i�j���wٹ��u�K�d��a�R t>��S��5V�{�#!V�V:_|�M%���B���>����*y�E��ȋ�)��6��~�J�;.�Ɔ�p+��u��Z%� &{"���?^FBȬ�6��Ʈ����i��Z��O���y�^�/��5��ޣ(��l����Ы+�lt���Y��nv�m��s�C46����5�6�Y��1���˫-S0�E��5+�A&��ݣ�1f�!]Ֆ[�W�R��2��е�c:Q��J�S�Y�q�i�mv�q�)�F9�Ԩ�͚@]�k�qdiM�����]����8(ECK\�d�-V�m�h�s�4�"-�;bi�ғkD��qe4A�%�5�n�@#i6�{��,`ZT��[IK[����.�+E���SfPØ:89	UԶ�@�B�B�K������t�9v'<�y��T;ܝ�Dj����Y�s�<�ml�ۃ�y��ϣ{|a���m�F�%�cGm��>���ճ []Q�U���!aI)w�����^#q0nw��~��5y����=߸��fs����8�0&2R�똱�ZZ	�lM�x������=uR��ÆG����	)EF��oZza=˗����{(��^_�ݳ���ͷ���h�]�7�������D��˧^%�^�Z��;�嫯 "p��@wz�a��i����SC�:�;�v:B]U^��,�5��0�[J��s>0�w#>���!
]��.�g���d�ٸѠ�
��T��b��9��G�7R�畿t�9�B�J���H��[v{N�Du����㞵��r�۞���93��Lⅾ���q7���p2�34��nzl\�� J���ި�x ѥ���g�K���������̙,�m�mnb19�M20�f�u�1�1;8��5}-��JImE�����%aH�ޓ����[X�U�ٺ��8
%���g�qM|h��p��̶�6��mCw.5n˘�p�X�{����M��6i(�Z��v����N��	K�����\��g�V��[�kG����Mw�5�bҭuj�����8���m��|��4Ǣ���zY�Du�S�y�@�Y��t��/��n酴���z���]�.�܉��'�\�ߊ�[3yx�N��Q�J(�M_���U;lßLd�E�����Ku������{��WW�0���A�i��)6ȚW��8�^"�om��t9�g����l���g�S��(׆_��������J��f��n�q~=�z�=��L�T8%��i�?{�d�平�9C��#ڡv�Y� �A>�{�g{�g� n��%f�b���3�8���$��ok_Rz����>��k��ϸ�U��"���<.���>%��{z2�V�#��q��3��®���5.h�47��b�h�g5����WW���7����{�m��j��+��)��"���i�ԱGEZ3Z�c���^�v6ȊDJА��C��laF�A%��7�Ҍ:��w��y�S9��O\��qЯO#���7k�ta�I!'���mk)���چ��P�}"���PÂ�I���'&]ٚ�<Ogu�\�a݌J�{�X�<kީ3��{��hӉ
�{�55�4(�3ܣ�"z��O�_R��i�sk���a�6��m���en�,Z}���"kd��s����#���W�.+�0 ��Q��ޢ��%���K��Nzg&�⍬����1⦕�Wl�F�KB�3:=�Ep�Z
�]Y=�k4�-�w���j���Q�V뷆Qt*�Z����=ֳ��Z<�H����b��|�Y%('���n&n'//Ps�{�&�W��o�z�9��tS�=�f�� 
�����H�:˕��OӺ���Po|�9�>��� �z��WP��JJ�`��G��
���)7d�i��y�HE#��=̝�
9�Dا�i�P���|�{Y�W֏�9�ˤ�i?Y��R��+��A̜��\0:�� �%��h�7K\�h�l�ң�0�,� �K�n�nb�e$��t��B,�uJ���>�wy���v�咝T��Ս�]�G�|�{T�`�$�{ޯ�����:O�ǹBQͫ�
^��)�
�i�6סMG e��lKs3?����KD�N�oݸ����ț��U�ы�&|��L�#x1���0:��m �L�Ny���LKgc�;�8��o5E�C)Bii��.��zu�cJ7�w�����C[	�-u۷S]
B������:;���svrbW��)�ZM]zd{78�]�G�Kִ�(ּ�ݹ%��R��)3ZEB��^�\iW�kR�	S���ʞ��莣Y��Q}��P= ɸ_y�;�����dm������`��@P�33�U����-3|��3n�5��gJ#�G�ߢ�<�sr��h�����5|2ga�򸷤�{��´eOlރ&7�,)������gY�H� ��/�+D�m��(&^R���㫻��U�5SL��ǐ�Q�w�����sXs�.�<��q��+��Ěp7��N3�e� eN8��G��U\b���=zоP�40���p�ĺ�B�@V�흦u�:�� ]�{�C�=�~������r7iy17�O�v�u�Tt�����ϝv�[��h�߸��S�93WQ@r	ݾ������|��eT��3s��f�hP��}�����G�'U�n�=aO�sF���ήf�Ou���v��xB�Us�kN{�����=~@,���PP�E�M8�
8���n�r��N^�=m��s��qB�u��3����������[�~pB���x��>ᮮHk"��Wz��q�A��@4��Z�;=]�_e��9�����u��z=�}ޗ�x��tǯ5�K�~�Lާ+niUOd?�d�щ�r��u��׊31N���o7���i��)�	!���c�+��sݞ�#��(�R 2_�%��A*ƶ��� b-7�R���_�z��7�J�vOy�LM;��������(���k��Tq&�❴�U3c����+Vj���i�yG/vݭq��8�<-�����Kǝb��Yi?��NRg(�'�&AS!Z��7׶���L-�V]�rƶe����ͬ�Ikm�9�b�P��ĸ��`+��(r�`Pؘ�M����1wV��4��e�m�x��B��u�lҚ�v�U���.�J��6�����Y�������Mj�j'	���+XW��k���
kiʆ�c�ұ�h�㭘)z\z�H��]ŻS:�[�T�tqeK�-S��ֽ���&��V��䮍��6Yn���6乀�6���sH�m�j8c���X����n��[������G���?%e]���F�qC�EL�5U���t�UK��f{�2OS�s�P{۷J�a�L�{z� �?({�P�@3K��4E��,~�DЅQ=�z{�t�D�M���ȸn�7�5����� $[|h׸��{����t"w�7�����]0�tĴ�Bn
�S~����E��ˋ>Tv��P���;B��N��"������F�j������{hQ�M6��l�^�>�[x.ڻ��%��*	�� �u7�:K�vjW��|w�i˜��D�q���#�B��`X5Z��[y�b�vc����ZU��'����*m�tΚ�5��l3� 2Z0�-���OP�(���=}�o�����;�=�q^1t�;z6��*�gOԎ	���V��|wث]s���J�W������ej��=����������-���Њi����1U���h
�ܒ�F#u]��,� [k�)(�	�{��}8�5=����wN��Ұ��xw�����4�֖��:r�k�gz���"��"zw�hq97韄���xup��M�e!���q��#��y;]n�9+$U�nzN�Ġ~Q��ȫ�5�nbn�;Ȍ���[��i������-�:͕r�D�pn�ѻ�/Н����s���t1������sƫ�^�9g�z�p��HM��B����s��Iŵ�^�w�9�!O]�PAr��|:&���j0�.=�;�8�_欘z�y:n�O�TM��Ζ焌!E�#6���w}>0�p���b]e{������d�#
�)��
y�5cbv��g�zA��ܭ��|�UǬ+Շ��>̊�ޯ�鮓R�w�x�J<}3E����Ln%�ɗr��b(M�j�D���w<z+A�ѻ��bx����dR-&P-�l�_�N(������qB\T��|ڟ;�̷�v��ս��U�d�JQ�us�1z�@�aE���KJ�n?�k�V���U�`�J�[�RXX:�\���6�F���{�).u]�1��4��F-��e0�e��:;!a����y���xq>�#@�&�$C{�n�U�Z��T;{Ϋ��ĸ⎹�C�'b�-Ƕ��2���ˠ�;W��hEl�D7%zlyrP!I:���/Y�h+�l\�{��������Í_`�캮�:{ZZcʇ����`����7��I �0d�U�jw�`Z�R�1�n����%�=�f�M�C(���S+'{i������_�ޟ���u���oD��;���%�p)��0��%)_�>��%�^:E�%N{�B��#�K���y~n�Ɨ,���s@��s�Lޖ�����q�AB�;kQ�� e�Q��[H���t�����e���Vh@V�`mX>Ĳv��ds���پ�q��2�or�#��km5f��=t`��^��XȺ��������4�N�M���=�p��!��\{Z�^Ӻ�wm�.��5hp�|�Ω�`�{ۉ�E�-�vɻ�.-��tU-��+����U|mh`�v�uKF�Vp2�е����\R���|VFv��f�.b�r�퍙X���Q]����
�۵5�Bv����N6z�$�a�ė3��h�h	�����vb�z���r-甮�;r���|�l��&bZ�K޻;�Ҹ�>��p�Xw��̻l:1�/��*�k� �E�k/N�I�u�lH��6� ;FuA�n�A����.G�.�3��	�-�̬ޱr�P7]۬d�4��H�^r����ts��� ���v�n�Ov
 Ԝgu-���Y�cY�Z�՜��}����Գ@�����}�D6d�s�:#��[�ybl"��\�3��}AJ=�?s���WS��M����	�x��[țޫ��8s�rۦ [�Ά�Ms�����ä���x�\�iu�:]ևz�LtW�S�F�Ay�vojNz=��˴*�ӧ����u��l�� �iuՀ.���{fŪ4�1��e:q�KYZw&j�7u���9�J�R���-�tdS�Vtɼ{��$(�d@�J���Q�nJ5E�'R���~�	Y��nh�x��K�� u>Ʀ�짣Yб����i"�p�I�ػ�G�|f�M����x<y��=�f�<��0;*_���*�_%F��F��U��yg���y���)z��/�݌O��[����B�(ܪ`BJY�����Zɾ̏F׹6M�ٿ	�r8ӯc���v;d&��g��Շi��JF	�=2�?[�sQލq����U]��F�9�5�=MW�J��m�Z�E�%��6����j@���k����Rm�lȗ�_OM���&�e6[s�l�'4���_`ȫ�*�B�ݾ5B�n�se�'^t�::�s�Fa��L�?0���y�SZ��De�='��pA#�aCKO����q���\�߸��+֎�Kj��� ���_Y��ެr�5x\��eK$�}(i6H���u��T�E�èy�g6������5G7��H�D���)�ïe��ǲ���=B(5�6&���FB�V���yÂ i��T�𘭵���5d�4��^�_�q�;��qvﰕ����i&ߍD���+Gc��b���ܖ�2���yg��� �#�e��3��7i߁q✊�sފ�#_~j0��s4�m�$;1y���ј�V�uxs*T��3)m�6�׳T�s#-G�����,�~�,�a7�y�ǐ39s�@���p��չ���p�"Ҹ�O��m�q[Qi����/K���g�ּ{��Ɠ�Ƹ��:z���S�5h�p��[~�7=1�.	�c��LQ|`�:�_��͌q6���+� ���֊۶�/�,���\��$��FYm�@�u���o #�������{;�,��������r�>�Q�]Y}��Ak^9ޅ-�\Q��zC/"���H؋`�}��׆x��{�_�b;�X@�%��5b��#l�J�|�©��w��H�"[��b���is0����o=��l\�b�DW>\c��ڡ�qg�6���/�z�-���׆�A��U�u�Gk�5�ӋMG-�~t!w&X5k�vy��퉎�'�3�n����{��һY������X����iCN֩��#�� [���r�\�X������}��p5���w�V�d9���yY��u.'��h�;U?�.�g��}F�*=�>��9���=�vn�M'}����
V�E��M��ʣ��Fu���rW;F&5)ysJ��+5��?z�z�j��w��Π�&�u}3hq��	+�v�,�]���[���<_
Yg��=5u�5!I�<m++Ԧ��\z�uGG{�(��;��=�w�|;����
j��������s�(	Õ!4�Jhy��	v0ځI�R�`-�\�غK��Y�雍y��)q����`Ħ��V�jLV�.YI��&#6�Ѱ��7;D�Ge��l��;du�p�j�ؐd�n�j�:PxG��Wv��è8ց�K.6�vb2�7:jɬ�\8��]e��rM�e�v�R%��ԯ,,2ꭆ-ѩ ������Z���(>_��\m��0[i
���je�ɪ�1�:�!l�q-����R��_-�aM�ѥ�Q%f�nv����˕�MnFai�����u���h�Kr)~��l��jzL���7�W����E�6�u��Tr�RO�S�1rzw�̧OkˬUVL�9��v�
���j�{~�}�n�rsx=EҁJ(�|草���{PfvJ���ռ��3��x�NFp���p���Rzh�J�_�2+����=*2��J:}�Dhq^�P3�k�����[_���vP��*+�E!V����]��	x2�=⧪��X���?xxv|2����7>���3�Ҿ��ċ�|:����~0KP�i$�2[VD�z\���5�8{0P<��g��|4��xW�����rn�+3����[�V����+�}Ѻ{����U/:aa�r�M�&�2I6)��3�
	=�N0�;w¦�	�2w#
�y�o ��s�O��uLp���hE�^M�����5�D-xė��u^U6�\^�{���dD��J4���6]�����Ȍt�ƌ��6�q��q����C�K��������♍Q.G=<�@=ڙ�"p�1����U�UO�F�����+�Ȃ�ծ�g�>N��{ט�{6
��,*3�z/&�d���n�l�ɱ�V%�q/}���7��_�gřC"Ԑ���֎�)[=��{�L
��S�Q�޾ڰ�afJWf��/j1&#|&)G�.��mX��]�}'�;�ؓ��%;&�1/Ϻ�$��>�͡[P�q/Pެ�^�sf�y��ѻ��{C>���HXe��i�Q��w��4Wm{��ۍ��7�^�j���7�:������F����� ��yp|���1�x�^�裱M��ez� ����6�7z�(�ݎ߰k�4f:������*q���[�1Q1�ɷ�*�%���h�g_`]�Z�bۖ�s]}��<\h�^���/Su""�9Q�W�Pd�]�hw�R�uc�r0�`˪Pqw�����d�Jm�p�q��cFy�O�MR6��U��#�(,��/�Yמ��]n���A�(���#��1l��.�W��[n�5��Z�V�,�N�$lm���B!�2�M���>���|�;�~�P2���;���{�R�^pc����_xJ*s�.O�Gb�4��s2��5�,fu����ui#	��V6HV:��ߌ�
И�׿|�?%�*5[���I.su�U7�L�),���pcH;2ϣ�O���*�̓�4���u�"����[�+f	���;����-(0�L��UC�8�]F�z3/�н;M�C���g���y�*��sǂ����?����ܾ��M�$�Kʗ݋jm=��2�K�]Yf�n��dJX�aZ����L�n��� �hթ�zs0UI�=)�9��O�55鷐LR�W��e�Z��F��f�B�N �d�M�"*����u�Z�6��z���f�F�����nީ�W��yCN�P�FIڞ�>�v'��k���y)â�n��t���P�-�j�\��}�\L�(�j�nf,n����P�_^O�Q�,j��K�u��1�D������Vv�I~"j��މ��8�-x��}��6{\H��7��]�5�ŀ��Ļ�T	��P��\h��%T��"���͖�#6�$�/����'Pn�W�謹�9������yM��b�t�?Z���Nb�/�R<&u�]G�^�^�/�+\��Rfτ£����O���M�t�R,�	��F��՞Oؒy����ƹ=W¡��%�9��Ш1�Q��>��j���V���3v ,��{:�"FlF�($	�y��@��i�{�����p!�N��g����"0H�/��j�:g	��F��\Vg��=��/�!h�*AY�K��8j)�T�*qo�GL(�-�Si�bcۼ�t.�˘�e�tɎ�����P>�,{2�M�q�5�o�:�z��t�a��+	�n�s�����*i�T�f���R���gj*N�5x��\�>_R˝וdI�Φ)��%n�I�;0h�c��Nl���KW>�1���ר���~E��� ��H�تDnYϰWήd���f�%;9�jF�1�b��5�OKs�@�t�}n�{/��"�C��	;S��(���#����ܩ�K�l�}�BP������������q�n���Xk4]iicq4r9�6u�BQ%!@���T~�/�}�,��w�40�_W�~�������/����Wx�A �����q��n��/P�]$8�� �Y��F���-���a�&��ooK���ѯK�����?�%�O�Go��d̋]�07ǧo�N�����	�m��IN�M�v
^X���F���E�nM���E�_g���ԃ�e�������|1��Չ��fsI��9_bE�f}[u<��!��LgWK����r_<��j���6�����7>�z^�K�e�V�����Ùxb/׭�W�4�G5�oƦ<�}�0lح/�� @~��"����}��}	1a��xg��4�PKM�%5Y��w�J���
;�q_Q��pf��s�q��ّ�txJ�P3or���2#}���ɛ�-�MpGM݁���	.T!p��8~[�yfv/O�"s�H�O�Yt4�B�ĩ�I�0~Y�Yx�E#���A�C�ẇb�n,ø*�X̸�N2��ɯ]h�!�V%f�#�K�5v��fv��5��b�na�ʋ2���L��{Ck�śD�,�M�2	��eՎ��\ivFd�J��^����U��.R[�$�K���e��	ihB�6�õ��F8?o�Bio�mteP�T�B%�aA#G.��sf�P��w)�[m��1xB�Vk����sR�F���2��@�Yf�&��9̨겮��5մ�hjn�id6�eɥ��ͭ����ݢR�ֈݵŔ5�R]�i�� ͠M��sm�4n�+aA��5-�V���c����S�~��s���	K f���3J�?��|`���~�>K��{kŻor�����-'�^h��/]����'�,�)���Z�{� o<���}���E���R����H�Y6gѥ��97�}�ӳf��b�ag��(�;=�	��g�y{���V�����S0&���B��$)h���R3��5"��UxO�Q�p��o�*Q���Y��3�J���>��K�.4�b$-���� bV�ʢ%��U�&l�g@+\mEdp�� ���������n5�|��K5͈��eM8L%�_���Gz��u%����w��b�g�rf.�����1�&б�]��y�b��)@�kY��=�S�Ƚ�{fP���+'��!ؽ�:�(yo�ޫ�VUI��+�7H�K��a�O��{��l3��L�ͦ��,��ʸ�VX�A�i��Z=����cY4�5����j.	G���
�ò@R�А���y�
�T�A�w��7R��\ӵc7������z$�:��Ή�O�5w�]�����ȉR���"�R�ICI�aA'����e!(�P���]��O�׼Ngc�/ ����-=m�0��/9��G��8λĴ:j��]�m��W�]�Gc���¸�^�c���r	�'b-`��� lv��5�V����2�n�.��Ϻ?��f��u���{�N��|�x?d�M.�|io�m�$"H�hH>���T�M�y����Ȏ�bt
��.3����6y-Y�媶:0���G5]�bwсY��F���캭$}�"-��C�g��$[LھW�ޒ>���~�O�;T����������^΅`f[��=+�������Y<8�}n�N��{w�{��r}Y8E�Ь&��m�݀�[���1��9������j�79Ƹ����Cbo	Ŵ�<���l@�Z���S�{�*lķφ��}]s���aqg35���-�V���?W���˥{%���V��6��v�v�6�]� ����.��ÝknI�ClkKKcgN#�b�a��]J��~�&�?C�{|��^�x����r6#��w'uoi�jt��.v�]c!XR$9���Ŷ�R�f��`U�|ݽ|�Ǿ�+�<)�U������G	9;s9���s�jGR�zԾR�V�%���%U�n���G-1|�7�9x��to��Te �,��x�ݷVN.��zПA����)�9���s��HM�-^���6�{4z'�W���V4g(�f_I{PfJ�⍴0�<��+9#a^=#�Y+�g;Uf,������O��]��4*��ƍS��_{ί��p/|�1սhfߖ��|Ӯ�3�9<�����u ~�rr�M�/���R�[^ �#R��o�у�}��OE3�9V���o��=��a] �ɕ3��<�AR�y��	��S۹�~���
�X�#f�U�"�^Ҝ�q�)��!s>�ĚB7��V�A�{���k;\Z�$�@�u�	3D`͘S�����Y~#c��8�b��XFjG++2����+])�i.���^�D����f����v�R��� ��y���WD��>Zs�U����?$�ʪgn�7���Y�}>��ۡ�5 �?��� ��UdcvT8(P1�M�K3�[��h��c������f*��wG�y�\�Z��K�?��7�\�{�:l!���H�Θ�F\���W�V!���Ty҂�C��Pi���T-��GP#ϭ�\�=1)�)�7���@6�3��}�8�XK�i�wf��{V^�������┺v��Za�W�GT!T4��{M�����:���{�f+��3�ا��fAVj�^|:j�&zqƍ~\4��ݡ[��U�q��{���+��B�|u�g�u�,=�+AA�;(��
] ��uM��:wu�RD��C"*�	\q�����J��{��4��t���HF�|�7	K�zub.	yFdx��SV14td�3сh^d�z�XU�;pD�A@p93�s}�Tu.3���v�n?�TScz�� �æS�E׊5}�yZ�=���Z��m�>n����[uI���$�Q[3]��j�����e�n�ɽ�
�G�ea�1�}��`ܘ}�:���y��:z�M������sJ�=*(�0r)
�蚜�Y^~
�g��H̙_.�h�{����ʆ�>q�!�H%��L7 �36�����>%�e	�����z{=��tʳ����M��kЋ�OED5p�*+�=�"��/�uyFgn�{m�33j.m�I�P�R�]�#c��rȾ��5�Ƙ�;8��~�T��$zf�lN�4�_�|���t!ufTg��G<Q�U��u��f矪�g�T����j&�D�6�p礉q�U��z.��{<=��u�)]̜+��������=.��V"�]<������u��G8����v����{��0`󷲭�-[�Q
�@)G�nkv�8A�;p�S��B;�0�����^�\a�M��l���ڭ��k��o�3J��OL�"�ecB*gz+��I����uV��c��:3h��%Rx��m�W7l"�����|묆ΜA�O��e�:L�64���~ŗD�j��9�2���Ks�lm��bѕw]��r����NM�����;�6�f}D�C����E]��(MA�Lߒ�L��X$���&�^�g��\6��|P�e]X�f���^-�C/']���Yu��`����-�W�rƍ��W���ݺ�g=8ξZ���c�y`.�)���ʛ�W�붥-�^�M�܀�1������G2�P���D+4�Y���V���l�sJpܗܗmJz����@���siů$40�pp)��e��ۘU.d�
z{��mJZ{W
���;��˕&@6w,�����P	:k.S�=Wce��A��˹�'l��0^��`�{�Y�r��k�Y�e���]�jǀ�l��@ԝ���F�w^�B��Q"�;#Բ�y�>R��W�tv���q;]2nV_k:���
�u�:�]�/�W��U��EN�pV���خ��lf��,!	`U��;�G2����e�v�>�I�8]0�]6�goG��"4���#�]Su�|���bǲ�-���A���z��kѕ/�]�f���*:���ˀ{���,�նh	3*�5�g���uZ�YeM��A/����vu�c:�sr��8�x�-n�cθ�<G��5��B%]D��&�f��͒�J�9YJ����avP�X�UF�����yu�Yew}[�,���F��ԶĶ���A���{c�D�B��3D����*o������ۻ��_G	{��ܳ���q��Q���ڭ8X���a[Mɴəh�.�ͣ^CR�ݪ��S1ų71��#����L�i@�vi�Ж�]K�C7׆;h��	L�Y��(7��kz陋6Z�vCK%2J����m�l�E���?M����i��6b�ٔ+5%���Ln,.�+en���Ъ��#f��l<J鮗M\鳥:�KH����m�c�d��ԥR�)��)�:Y� �����K���iY��k��� -�c4 �p�Y4�6��ˮ�K��ږj���٭�Ļ��F�v�4� ��ԡc��it�;S%cZ�M�˃[[x&Y�������B���ҬSYL�Fk�����v4Wbᶱ�Jk��cMk!*h��j����u�V�Z76��
H[Zகڳͭ�9���#�:�d����g[LjTع �6�-�����W"V��f�Y	vu���$��YCfۭ�]z�,tE,-u �RYL$E"�/!]U���C.6��ɶ.�XK-e%Ŗ�.ڑ	-�KBm6�*#S:ZV�af����`�
M��2�yiͻ�Jhc<�ViucNv*D&v�bR�)vָ[pn`aF�ˁc5��jJ��e�ۥK)I���eͅŹ�f�6�h�M�P��G	�WZbf�.�RV�+-�kf�j���6)��.�����-�v%��b`rб�*ɶU�E�����+F%ŕ53%G�a�l4��	�V�9P�֖�^�À"�n,;׭Ϻ���:�G/TD�Ԏ���S;1l�jBV��3�`�iȡZ]�PУ6���:��`��V�Ҳ���̻YH����Q�c�[d���I�-�V�#ce��0�� #�6�Զ]����ӈ�8����&�a���,]�Qu��c�\����f5�.��_y�]�A�m�C]�(�a�{@��2�vy�L�ul*˃\[���&�R���&ո�ٵٵ�/1�f�����W7&m�����#s
MӁ�لy�]�q��ˣpg\SWV`L�(�T��Ch�(]s��vfe����2�m�ц�Xe�8���v���rVa��l#��4U۵���ޱ�\��ɓ5� \L�فnB[i��l���e�.�shl޵@�b�,��1�:h��^�j�һc�usuX�]�)R��&�Y.��bRVgYn��*aԕb�{7]F`{Jf�ҊCQ�6�Q��i��)l��x�ީ m�l�78	5�ii�[-�	V�b�	��g,�tu��"�X0�B]h��70��M�����2��5R��*5�M4#�,5��&�cd�;[e���I]u�u�h�f���ˡ5���Y��̵%r���M�	2i�8�\����;G#��122����I�M.>�)�����*co��UFΟ���da����oݕ m�p�uּ(g`�2P����"�eO���OW-_lS��<�g�A�5�L�{��*C5�}y$�3�� v�\��n:L��D�8x ��Һ�����.�*��_/V)�q���6V�F�\���|�r����	CI˴O}�L��A1��	�#��Ȝ����kK���Q�	O�v�E��sG�6oZ���i�3�p���&U@r�N+���Bgt�W,=�$"���S���:J�Ն��.S��T��Mcc��׹L��n`��`w��N��6��U<�.����Ĥ�L�s����P� 8-�Si�qbϼ�l�,x���5'��3FO���[/ϵ�j�\�����# !K���y�5O�4Z�z$TU�w;�'ِ�TgF^�WN@�h��3cd&�]]@&��ģf���)��n��ܙؤ\�4]�UH���"Ȅ"*VU`7��_*�5-�4΅�y#s3L�J��[)ל٩�놈dހ�=�>���7��Nd-�-�����O�Uό�n��%��?D:�d��RP��ɒC���yV}��=��<M#�_��ea���|�L]��o4
���,%]9yQ:�#MZ�T��2)�\����Z)cB����5�9�X�ѻ�̌�.�_wRᛙ���B��}��$�Z����o.'l��v{j�|��K���--<Wk��^�w%tt�j�XU@1����'d�v\^Iu �¶�6��U�)�~�Y蕱@D�dH�\�g�ը��2��Ӿ�6>�V��;�:��=T��9)Ck{���иs����V�]����.lL^�l�ڟD�:�?UdWjc��{���td�8��ڼ��0إ3�4���z�ou�;Ʒ�;&��E),$'2-�߻�{+8�7�g�R� �����eow+�B`����,���S�3��6&q0l������U?G�Q�2���q���i��e�i�%�5��*Rh��0%�r��4Gv�m8��莊�<Cv�<�~�F*���h�]uG�&�v��z=���Gi�b���h��q����ԮĨ��9��"�"p�"�o2�w�a>�����Ua��zc��e�{��e�Ƅ�g�Y������w��1_T�tI��*!,�e?��Tᰓ���)��g/g�s�+�:�f�7�zG�c��3��td�b�$��Z=�J�f���m�r���rc+�Ux�
/�.Ř��Y�K'
}���gt}ֈԠ�V�V���j�7�ʲ��b�E(5�
�l�7���KE2X(��(N��3;<n�fWK<S�x�C/�����ݝπ�H�t�]���ko���?o� �3�k=�>��t�me�e�!\�ÝA�&	��M��^
��~����^�ɏF�wo�{�Sڌ�3��U�o"zW����.0�����uL���zY�N	��(��j�(�����g�%���!�+-�ui	�]K�l���\#R�'V�4�ȷ���w�ӳ^��h�וJ�L.��7�yeb�.�$o���GW��O�X��ެ/V�H4K
�h]ַ�A�]�*��b��:����f����B������{��旙�=i{Wm���/]�:v*Ƌ�7�n������N��D�H�f�yߠl��h_tN
�O���n$��ꑳ��Z��4w�z8S��u���_�\�ޏ_��5ӚK��&����`�A,�*�\�OGT-^2�������3���뜓Qu�LŽ]�F���d���;g3X�Ӄ�B��ͫw\z�_fԡ\B�}g�h��N�\kv�4p��y�f*��V�A�M���2C�U�!�,�yL��/�uӫ\9N���:�fLn�Ρ���}��M&}h�
@�-�����*X���[9q,`�����/�X�ꙣ�s�`�U,�|%V��ɿ�_[t�d�ܟ}"W��g�=Mh8��n�,�$�m��l��Sf�ʐfѻZ8(�r7`�
�[+��C�\�s�/�w�ft��>���}T=��z�9��&V�W�H���
}��tƃv�yw��ٮ�X2��C��3���|$ƨ��l�Ç�2SH�܆����f��M|�}ǧ�7ޤ��K��ޱ2<��"b�{����X�[
l�ӂ�4[U����d�V�]}�2T{Pu�}>�:��]`љ����+�ۺ{�6Zn��6��R���L���U�Y�^c�	�"`WZ��؜��	5��8��V�u�ck�yxh�x���=�U�|�:�UBX�t���
�++</�1M�{�}��y�0�hA@����}��ozf�5/cM�	��Q�Nc�v���H��y��w���#ڽ��t��y��j_���������<�e���Y����K*b����{s+3N�h��MN���Ι�zٱ����2J�Ĕ�˻eoU�ܗj�oi?���"εߜ�Ҽ�Z�n�X�Q(�u��J'����4��Q�`n��vҁ-vElt�$GWmCMnnIw6�ڱ%��V��͊J���km�l����*��Ys,f�v���1�ݶR���0Kc�]5ʕ���
�B¸��v!Zv���XbZ�m������6���R�@Ɣ��Fj���a���L?g�{Ε�I�CD�kؘ���WV*�m)WQs�)���.�AMnƌts4�-r.YtƠ�[LRE,WZ��Sm�t&`CZ��.��3����cS�M:��r���ɖ��X����R��@��<�{���1¿9�T�d^:�˸;���:��������gX@�b#��  ��G��K���n~Cl#�\4.�WQرFfz����c���x���3� ���~r��T��A.���!�	pY��w�nzܩn��Du��{������Wٵ.��8@��x���?g�i�/��ױF��1�l�&��ϸhs��ɟ%n��Ӈti�j�yF��,�7=ߺ��U<���.ܼ��<��0��vr���N����=L(h[��L�����痎�Gm[�����.S�|��9�`H�#j�>��v��n@���gT򞧡�|)�P+��t6�T��2���&�kl[M�YI�Vl�!�M5vZkur�tQ��oW��+�wԫ��䱑�V��]VF�6�_zٜ�]�FNmUȒ��S7^���8߸����"B�-(��@�;��l��	��͢�v�1]�@g���px2©��)\ћ.��
ߴ{���%���Yf�{�����ïue�����������د��Ev˜�o���;�p�΍q������tx��I^�U�o<�ȭ^��:ʼ��FL{B	��P����Yk���=1�>K��z�Z�}P�6���t�{pt��r4� �V�ջ=�z�ڟes�=�F�h�� $���f��������ゼٚ�
�؂����r��O�e�w\�s��~���v
�"��O�	��
�޻�*Њ*��w{ֽq��:y����~�>�x��%t,O�QO���*�#J�ԏ<2=�����ײ%w3�ޣ��k64^�\��5k��q6�T#�3lH\f�Ҥrv6�̚t�n���h�����2���br��Ǉ��4'����{�949��]L��c�U�
W��8�Ig,x�ε��{�Xܘ�ja�H�E6��Ƕ���ɮ5�I�}�f���;S9���ޘ~��˱�n���jC�����w�ZqƮ�䨒��>&����㌬v�4��"���ǰoNE���Lu��\��U�ygG�ǳN(q{2;�k4�W�ꑨ� [(��^�g@���Xc@���i��x>f�J8�9��\��1<=һ�43ݷ�ky�$�!q���l���_��^����Ϧ=����9��qNʴ)p@�Dt�9����<�G��R�>O��O��,��w{�=f-���z��s���=�Z�1�}�׫B�/?��P)/&d�2Ji��OJ������G�e������9������1�W[ʔV�8E	�ڎY|��0!�B�,�2�VN�E��B�e�º�TVH5`��ڻF��kY�!���l�b.DĪ���Աu\��2HP=�֋���9�����^x����
��W^v�U*9��*�}��k|��Q~����"Sg��{;���ǞnJ���{-6JM��	���&�n�=�'�Ȏ����f��S�b^�L�Ns��T�mR˝<���[�B�[UKwk�4ԮFV�R�.|��hɾ�w��O����7�}w�ʀm�Q{��\�o��*6o�̓��ڙ[� �7 +]%�5�c3��� ���5��}y�J���%��%�~��a
�W�w��v����OZ�H���ۃ~^���U1e�1ߔ�6j���c�8#1K9o�e���
VnJ���	b���ZS���v9|�*���NV.{�(�$�2��^fR���ِT�l5	�*[��U������^/\�
��g%�A�Yާ��Pi�Ȟ��Ќ�]��*2��pg�v?:rH����h4�P�N0j@�(��K����A)�6�	����骍�����F!:Vϊ6�I���}�����z=�؟(�<��x�p�*���S�`���K1�zc�]8t�1GF�H���Q@6 �M���i_V{�f:�}KX�!���tMD��ى��7�n�:�\��ES�#W���G����;z�t
ɾ���i��CNd�(,�(��uXPr��y�|�r�r9���򖬸��j�"���}�����a����K�͐��U҈��#c�4J���FI�Q�K�eȦTӋ���)��ֲh���?^�,D��۞���~���(S�{b7+n�����p�4����-�,8A6j�=>����v����7�������M�>����k��� ��l����'O������/G?�ې��ʷ~Ϯ����&��9})���sD��In�weu'4n�L�q՜̵s�3C�n��+��e꾘U�X��3�l�d��M�m���\�[k�v���؃�*8�j�Q�Ken��Ĭ\h��f*M\-�ʹ%�(ʺj�^sZڶ\4Ų�0��kc�C�%�ݫ.����D�NYm5�֖����[�@j�h]�m�U�V�lX��-�5��αv��h��̩��d��7�YrjJ��p�"K�f;5̨fg)s�3�)�`04�^�ۭ����+[n�]��vͅ7_��؋2��غ�e����W%�����2�,u�7A���KU
\M��1h�s*[�A�t�L&�d�������s1���ۊl��~��t��M*�N�>�W��0pmM䂮��Tm���~�e�����{K#���"���G��YE���Y���<@v���f�&g��Y��΋�����F�vo�Y7o�`�%��2�oe��n8bp
WT��t��h�5A����9(G��A�0,����[��#�ã�~�Pf���8�(���϶��9�w~Y��Q�g��Ǎ�.Vȉ.��l<�5O����p[�缪�lU\)�+Ww��NSѸ/x���70�P��n�b���S�<'}�5#p["+b�@�p���޸��\}��u����r}s7DT��^�w}ũ��&���|#�s7�s�W��/qz(\2*��ڑ�k�0��WA3G��/^�����k�X�"a,,�	U���T�>����z�m��{���uI�k�6O6z��:"�+d=��h�����x��x}�j�>�y��d�:�X�\_k
{Qv��]����fM��S���g����P뮣c��AUpYt(�
�3X�RYؒͧ��+f��繷A�>33��,7u,������(u��epf\N�J����f��N�y��^�Q�||}��?gd�=	�+�<�D��w���f)d�&�fW�=�2+��tjZ�͡q�>DToݰ�U���Ŷ�&�F:<7g�����m�/���P�ie2!0�M��\c��]�����r\ޡw7+@��}�vw�<�}���H����/���7g-�mx̫	T�Դ� K_&���DO�.΃}��~��i� g �rdml�9�/�Uynm���l�v��Z�N����\�\�tK�;10Y Bn�
�YTk�A�icV��ڹ�6�ͅ�nm���kMli�[��~��3����>�x��8����s��mv닋G��2�s�#�f'dl�Ȱa'�o��A�=8�LgT]ӄ@L"�)��L��\S�A�z��r/7o�l9{T�U��s�#~>�WUv�����~>�~46+�����}���@��P�M6��l]���z����X���V2Η���r���S���&�������P����г6��.B�张�fjs~P�MN�9Fj/c���fTjt\��s�s$�������q+��~ݫ��A9�'[y^
ξ�H��,>�Et�ub�o��x�m�|�(�ޫ�*�߯U��wX;N63FJ`���h���c�Ҥ�͟�A6�mv�R�ǁ%Қ���J�槀	j����:m����m=�������Khq���k&RA��=1��i@6��l�B
���\�{U���y��{<�2�-B��b��8fAi^�a�Hʳ3��w�UիS�ɣ�� ��C`ǒrQZC����aD���w^7�1fɈ�K���;�����V��u�����═qRg�{�`�tq\�ͬf�l�K��P�:�D:�{A�R�>5xpb�|�/����u��+kn��y[WWpVRC�\�N��l9�I	��4��拮�4)�PL��휬=V��ٕ�#��g��b�gq۽��C���%�|��f��iV��U�3�d��3����:�v�KV[&����f�Y����
�1��s�W`��n#d��殃�j���(��:��/5����RQ2�+�-R*Iky��ۗ��ĝO���V����L����R�j�1�y�s3B�5R���W���]�`+�����xT84 �%�[�����1#G&ew[o�w�)��76��7c׻��Lp�;1w@�P
@��d�t���M�TC5��kbV朄���]�EY]�\̌�kA���z�k��V�pe� eZ�Y��F�J��6�曆s�+:R\�+��W���K+jS���y"��
��m��lgL�5�-ž�[w��\��Y�d !�p�d�]�oתM���o�_@�dy����3*��"e�1o��ZL�=:Xu���ґ��Lt��o�3��^������e�T�Lnk��4�����E8�7���V��O?Z����{θ-~k�Xo�χ>�x�ce��d�Z�x̩�+�Tҹ�%���[�[W��s/m��f6�bJX1�����_�t�����7h.�?}�9����V��1�����{�rc�������=��;ƣ&�7]�e{i��Y8>⓯;z߶���-ce ��i�~�Xs���d?:R���[I���)<�Ә�g&�7TS���LV��NOC��'Exk���9Fܚrr�aD�@$6�A4�5�4�;v��fh���������!��|6�w���S����v��ݝp���9Ex�]BV.���è�����+VW��b�y�R��RsY��#޹�k/��ז2��C����_ݿ�h����� �j���G"yn-�'ڜ;)A����jq7�-Lb����̡{�Wn^#�PI��ot�3�燫���	����~���g_�BBL1F!�VRGiA믷�C�ú��;|;X�������|]��z+��d�ۡ*=�_�1���Zk�\;����/=�Z�yw�Ztp��N��7�=���Xf� �/F1j�F�Ґ�r���Q�6j&Km�l�����Ӣ�^ޱ������!C{���~�'�E�j����"ɦ�;ˏAο#�t�n=���x�6 (M�k�(H��`��7�R�̈s�4>�xF����טb��_��nr��0��Tnc`d�9C��f�؝���S�r��+��r���UUT��Evl_SaU��&j����5D�_{���K��7�9W��$au6�b��!��� H���yO]�I�ni�l���
w'޻>b1ml/d�s{�o<�E����Y�Z���jj��hk���.SKy���x����� ���_y��CI��m�]��S�xJ��tUĿ���-���G�UMZ��΢}#Nʞ�m��:�z��α7?{}0{uר�?l�>X�Y�vKn�[�3E_���C&\	^3o�̓阗������n1��^�"3i��:��-�C1\v�<��8s�ø�&/��.�qEQKcc-�T�Ѳݩ�t�-�Қ�u��\Y�6Լk��[mĵ
T�Ym5t����E�g.��f�]��nS\��r�G`���eu����%��F�h��[.�j�Na�S-�݌%�b����[4�9��ln�kl�Vђ�k.�n����a���E\�KsVk����Lnnk^�����1��fs�چ�a�n��d���������j��M��7bP�����.�0�4���Ԍ�t�Ĩܸ�l`�Jf��3�eF�[�Ͻ�S;P�	n��~Ϗ�{.afs�?\�l�������U���v��Xs"�6W�����������ݨ��y���l�>
��c��ޜ�TV�G=B��|er����Lfn�}뉾p�A��B3^S,�w�w�D�{g+lC�Ņ�+��,%?��i��3�}i�ֱ�1[��8���1K�%O�[y�2A�@�+�F������f\�N�0��QU=�}Q�,F֬�W�!�)��G ��������*�х�X7��U��.�nxh��C:g#}�}�aw��?w�[3�=y3p����)Q}"����/�}�n��(G�	$�k������>���g{n��Rwo����۝���˼2=�^��9U�Da�%uAwe{w���oq<�Q�} ������o�����\٦P�c�6��%��Kn�/\/G[�/T���Ɩ 1R\����&u��C��>�{�Vw%�پSc{ٝ�r�-Z�O�mZ�2uc��U'�S�������� � }�����`E�SD���e��#�{{��݇�6g����?�P��pyЩ�Q͖�nKb��'٘�1p.̨uӳ�e
�ty6"���Dmf�� fY8�up�~�s�*�p�lV��7"}�,�e,��W����@��=,ҍ�S��������7�sl��i􎈎t����{'+����=.	���Mwa�R�6+3�!E*ܚ;qCv�ʯ���~���l.���B����!JD�(7}�����,���R��G��uxOMD�V�aL{ҙZLyox�ڃo����+�Yny�E�k�W�^g��V�{�.=1��*
�Y�h��U���5|w���Ez����]�W�N���; �h���z_خ�-۩Οw���z�S�'��z��O��g�{��FnL�ά����&jdlt&�f��@5e����L��j�7��3���R�L��I6}�YU��T_�\Ѿn���w6�b���^�IwkgkH{אS�nW���1��#��_��颣B�Z!�2t���(�\
;��ޞ��;��v!H1u�3�
�v8̌ǹ���qt�;�E�x�~�����a/����"�);���SnG�EJ�������U���=�V-Z\�����̉~�n�~���YC�iI�+*m{{�co4,�,Y��-�J3�����{Y����
y+�ey�g�c��7����Lף�� �gpW��=�����^ݕl���ޝ^����Պ�1�)W �o�7 �Gm�)�ډ��cb���h�]�h������ɣ�?����7�F�g���oo�w��O�P���)�X��ǰR�/�r��2D7�Kv�%�s�V^��C�}�; N�V\M��{�(Ul*�s�&E�M����"���e�K���:�^ل�C32���-��Q/���k�Uej�U�����P/WT�5��mk}�1��
��S���u{�TPzgZ�.��Y����n�=�3�Q�����\9q��LJ�$>�
��:��{���չ<��aWLߦ�C�؊�n��}��$�mZ��Cg�?�[z��2+��s�$��%>^ܛ.�:IH�4�ls��r��7t8p:�/+��n$fd���Lg?G�<�F��}ˣ�Uvٟq4r���{���S��~\RÂ�l�v�եN����dy��6�;�off	��C~�$�����d�-5oW����vɭ����q�"�B94ч��NO���j�x�����b�F$kD�d0w7���������s�	�t�+���-uO�"A�_V����T�m����> ��N���b��pv-2������[�G���[|��ݸ\۪~&�:��cgs�u��oU��z�Q|���G��^V���t��3X��U4B5A>��..��0qoU�.���+t{`̠�D�3��iq��b���3�X���{�7�c�4E�������O����/:v(ƺ��t��9W��ь����	�-���}q��l��?Tu�5��%w~B��V�������2k¥CCϩ�8|�5��=�'�ǖfWEL�D�����
�ߤ�j2�Y��+=wqOg�"�Kށ=�~��}oc�.�y!��v���l�s���M���:����/ХR{iF���![%�5z/���YNJ}�]��V�}[j�_�k���O{�N��;goqG�Yo�v}���*��̺K���W�0�ދu����	m�\!)��=��"��CO;����,�0������}���VTZ)��)����֙�7�~�hs�z�����iS�%�^B�b�=���$=y���1��hu�էdf�_gX�:�F,Q�-3��[�F��M1�Xfں-�e%RQ�:�$h�
|�,\�]-��5���%�vi����m�w�hY���+%�!y�V�Ĺ����cy8�Cb�\�����Yd��<�'U�=i6�c0[�R�$v�N��)x�b��蒥�\<u��G+*ŵ��0�t�;C)�v�=�#�4u��5��XM�5�	q/,�/>���B�Ĕ"�)t��WGZ4a�\����52cl��esY�UR68q�%R͍ؐ�S�0����²�A�æ�Y�r6����ިB����1Y��"ޥ�kB�5��	���X��f����g��W�������(�򎌲e��(i4BM���MvH���7ST\�q����~��x<2&맯�>�N�\J���ԧK���P4��2;ѷѭ��c��h��6�&����GV omOT�����W�vjg����p}+I�cz��3*i��C��g��Z*Xfp[	��i�ޔ�H�b�*�}Rj�m�1�x�Ψ��zb�qIlN�>�~�w�Q{S�\u_�R�]Hi0�Իx�:��#�_n��")��,��,t��ڏng+u��4�{�:�*�:�)�{����+�����kzz����Mk�bN��~]]��]la�G�]�B�*:�Kљ�Z�j�J�L��7	��7O��2�H�O�e�/�>pTa}�����>��|��x#W�w�[S�67@a�~�Ɔu_8^��S�G(�>f:4� ��m2ٍ�������T��^`���f�j(k�Z�T���ye���i뎧n���s����m���ޣtf1;\㠋�z3��(����7��U�{���U�^�V%5��	���;�B�_`v}[��᫫7��e�{�LO[ћʱ�,��)7ǫ�?groo���,h���T�GE���A�g���i�×�����}�7s�u�����W>D2�0 &��o�N�]		u;wfի����z&�Ws�y��utkGY��[2�aɯd��]���ʀ����S	(	���%�wj4��[�Ƽ�G{ȉط��+n
�3��®�ϮU�Z�T���k"��'b�d_]��яe����Z�ĥ�$�SH�u��Vh�t5S���۵.[K�۰L���n���M�����1�T�OO\��k�sQ��}�Au�s���v�g�[�h8�"�6��me�l�����	����b�yaQFD�l����]���v�����Z{��^��ˤ+�M��-T*�_*<6�̸�㴩_���V�Fvݟ��
�� J?�i�;�X�}[WԶ/�|���D^��/R=���y#�_�־xA�|m:��r���b����Ƭա}�{�%;�F$� �Z����[U�L���b����);�6�oL�գk���Q�[��f�D]6��_� Ԯ�|��)�0ᆜm�J���z%�ޗ��m��́ȹ����5�}v����Tp��T��hƺeZ��9c%�Sv�
Q�Y���a�nl��p�I��p��9��q&���U"V*v�E����\�a��W_T��OFӗ�_)��R��nv���|��7�"-y�ދ�i�o�#�B#�P�H�i�iI�0u��F�6��GU�q���\
;me��F� ,6��~y�ΕlzWi�z���^��^��v��%g�Y����y�R��+�w\��C
�;�>6e��H6!2Ym'گ��S8n}��Μ��7qLY�upH��ḱ]����?U�lu_�P�|��z/p���d�8IY�6�\\�����qB���h��=@�rMf6���>��c��U>�?)���B�7����CK}S���o:s�n!��z}ȫȝ�{��[�B
�(� ��^�+�3�*ZJ̩�~'��%l�J�t����Ov\=���n3��/�w��q�þV�B/��:�e�h��x�S'r�q���e�g�b�Inw뵧�7�vr�d�^t�&�G����;�Co�MH�L�/۱�=o�u��?���?�2�Y�F���/���k��u�����D��uәQ��U��3���m�w1������\�����`�s���R�����bu���vܥ��[�n^�*��eK5��M�]kl����SR�ݑ�v��[B���sa=_z*x�}rf�ش�8����cxVe6,�yVy�[����
c����r�&l�F4�pAm$�-5谪W��ğk�]J������k`�Sr-����s��]����=؜��pvX�Ls���}�\I��խ��=�w}Lb �
Z���������Ү}.[��1C$��>껎5�5��\	�Q3Q�}��.'�E�׵J����2�Tve�q�]�iHI ÀXE�%��Ye��;�3���G��|�����I�u]�N��-��C{bwE�Ua�R@�����ۛ����پ�jX�K RKX�i�|������������̋���9�-��I���$��'2L�I�m�k�۱{cY-�m��7��v/!EAW��APU����zQs� ��H((#����2AEB�
�䂀 g� b"���c��(*
�g]�8�WG�֞���׼�f�yn�Tq�u�c�>����"*
�!�y��G��N�����k����DT|:�mҺ�!_R>��f�����O/�����F���ןL��E�H ��h"�	@Ȥ�Ȓ/�%R) 2"������
�
�H*�U��} ���"��*�� .@E�
*����H��$��  2*$� ��H�"�0��� ��"$�� ��(� ��H"H�"�Ȥ�2(�2�H��HȒ�"�# HH���"�H��2!v�(}?0EAW��Z���������/]�sw�O���M�y"*
��W-֒���O��ӕ��=�x���Ç��_Q��8zA^'0���Z?�Nà��**
�_G�p�l� ����9k��4U�/ꈊ��!_�%����'�s���9Bm����n�������rQ� ���>z!�����&��������������*�m���	���*�=��x���56x[B�qjӶm|���/o��(�N��*
��|%[���`Z�]:rg��'o-6�lc��PU��b��<:z<��A^Ӂ��^�v��;:v��;�\�����)��1 e��9,����������1'}��)E R R��J"*�(*�I)!"E($�(�J
����U ��� �E$TR$����J�$�q� ( �  �               P  �((       ��RZRJ�i&�
Z�R�P������
��*R�J�R���� V� *��(��D�
@  
 P ( ��d��^s.Vhi�!�ª��Ԋ�eɮٖEe� �M�1�j��9:�D6���u&�{�z�f� .핚��wk-�ͷ,�6  � � �  �����=�����B���
(P��:<A��(x� k�C�  z-��� t^��5�myܸf����깉�ڜv+���6:-�� � �q�PA@   P w�Q$�4�F����6�l�-(�Z�]�c��9UW-�Ʈ�͋�8���Z�9�f�5��R��\ c�l�����bW=�hh  �����Tm����-���uI�:y��+o=�Q�2[yt����.6�eQ�p�{���Ukw��,�N-�d���
3��E*04P PR�@  @  U ={j��nز$�=�W��i�w��	d˖�d�p�{���֧{��l�֬l�W.T]���.@�Af�:��\�9m��k���T� q��˻l����J� �Uu�r�՘\���j�ȫ���w�Y���(�U{��Rh9r���)��R���yh�.̀ B� � B�   ��iM���m��s�lӋ�m��ܺr6�iǠ�/l������Rۓ��&Y�:���.歶�˞��{j�ܺ��)K�˰  m��wjR�K�95�� ��KmNZ��'�f��������l$���ν����r;JM�ݚb[m�t�LTrݪR��@
�  �@  ��y[i.s8�J9����x��4R�8��8� 1�@R����s)NZ\�A�E����Z˻V�y��^% )j�4�y�@y�� x�Fv z�s��fµ�Ɣ�#c���@f� p4
3��04��^��� �c��ϩ  @ �@jR�@       E?!�)RP�0&� L!�0)" Mid�h&CF�M�FԄOb�H�I@!� �&�a0��� �?&�T��0 L     	OD�MR��z�@ hd2  w����l�yyz��9��͗>;�?=iѮ��m�:5���
��u�1�;�;�٘`fa�O:	ç6�����xɅ�-�"�2J�/Ã1�e�D��)P���������/��_�ݦ���S�fe�Hܕ)Y4��K�4��]y+eb[�2���33a���"�rͱz�Sß�gc����������ݜ�n\�IR��X����]�rh��߅���z����z��L�oy8  0���������5�$�����=��뗕�jY��8��Lf�ޭ)��7�
ٓ"b|��M^��ܠ��2L��4]ia�1�Pfm
E����w���i�M�Z��p��fJY��햱� �F��貞�˽����0e�1Zj��h%Q��طy6=���Li�������G[�LѰ�3fëfH��ђ�k(����(�xN:���y)A���
�X�k�"UH��iWt1ީj�W@i��m�`�ŖNѡ��&���)��!��ؼa5X�M����B�m*��ܦ4�;�R�u.��8ּێބ�n6�0�i�oٹ(+
���m]D�-mP�yL�ŵ����kb7zS��6�IV-�-P��!�k4H�ʻ�5ѩ/j��;�	&L�סO�#b������
�Uu�2`��#wF�<yQh�ǥS`<��ˑ+�u�2^����'�����F�G�t��j�V�ZZd St�T&Tcof��J�`���j��!�N��{�̦K��l�x;����4�Tb���m��\��m���P�Y-�UôC�!R�|i�e�n�PE2��x���*�V�f�Q��{oZw^9NS�̡T��^���baD��L��ض���r��V^���u!��^՛
��B�<��%�S�5a�A�d��ZQ�N�̻OT�E���Q��l��h:��#r�L�b��H��0�M8i�s4L͛��	5OF��X���pJwq�v�K �Y�p7�Zd��v@gE���up��
h+�B�cL7��SaZ&�JU��M���bx%
��֬����e�Nˊ��7>��2M�oi�ct����y[�Ѧ�\2�5,VU]ղ�;I�II-�ǖ�m�3&F�� �;n��=�ec�+$�zQm*p['n�㸃ە�M�"�N͵p�`nW��� �e:�r	��97Z�I����*�������2�@���*
�Wi�A:њ��+4�Il�;�᷊�d�n�m�-5Z�5:_]⊲��l�t���j����[��v�� �����:��N�Ur������w�][�[��* ���u{phq5K%�˵/����cP��i�ͽ�Aw7d���ǳF�]"L�.��Є��+ihHҫe�)9D�Y���I)��YTc�R�P�U-}�(Ǘb�Ѻ�)H�X���Ѻ :X�5�WX1���!�[w�8,(%�kV�kV�Y�fm�EJ��<x.�n�C���!KJ����8����  ��9qkv�x�<ZȰ��qDL�w�7���cØ���q�B�8�����9�Gk76nˢo���J�YH�Cj��C=�6	��f%S"�0��ljJ�h*U��2�%���գ[������D�L+d���&�7z5-�P���dB��
��c"���^�6!�����U�x�۸MW3� �;)Tc�I3�ڱ�Pgo�Y�dB�3�m5�Iݪ�*���t��fF�,$7om��ګ]V��;�vʖ��`v3H�h���KpW:"�,Q9�%����D��ش�&�cE8R�,�M�)aZ-��cZה�'i�"���Ee�\��+f��i�<J�[p[!�ۦk7^9@�S�QUZ��
��$Փ*¸w9�[Ҧf��v��i�{�ZV;#,�ē'��SIL�ܔ��*��"�+��] ^�{��ZB��,�1w�l'�ma)��(��ֽs�5 �V�L�{��aQ�mw�0m��7{�kh�+u�6��-��`�^���	nU�*�V�˨���j�ר�����q��n��IZİ��Z��8~�S6���Z]�{A��C&Ņ/]5-���B����/����V�@$��u,\b ��r��vnwK^ x����fJ�X1���n�-�	iv쳑ք�.��"��eb���S�`QKJt�76�ɷH�3�>�Y�P�+,bێͷ�~��m#LbJ��/���5�Xj�H)��֕4Hiȶ�P�;D-*�F���Y�)��.n�t�%��>��z	��	��j����636Ky@���K��wqJ�����gHU�;kreɑ\�V���E�5Ԙ���5���/E�t�u��X�V�v\�s%VJyM̖1V�u�hC���6�B�Ԃ���V�aQ�\�Gj�-J6u��x�w�:���bB(%Pڙx�ya��w7e7t��2d�N�������r���3Vj��fmʼ)��z
#X%9Xr&�E=�z�j���b���[��]j�j�Z2��*k*�5ۨꢪ��xr�F-�(\-��3nV�������A�R7��`�B�[X2ܩ�."uvӷ�F
��Ytr��h���ڻ֞�Ym|U�'wcѭG��������GQ��H���rլ���(�b[�cH�A����s2���6�Qs,݌V`܂���t��z+Dk�ʘ�����ێ V^ʲ�pj,�&��Wf�,z�1:�M*K'R�h�W��4��mǏ#��$Y�U'X��^�iɛj�ōK��3���X��6S�s-�`]8,a�7b+�j�Ī�x�C�w$�^
��Kz���o"���H��6U��br�:5]�9e]m�vR��R�@l�D��jX�,�G	�(��٣K>b�Ew���ނ/�"!hTq�ȭ�9D����!��iù��;rY[j�&P�l2��)Ud.�Smb�0�̲^h���@�ZBѩDL��^�a�F���tMY
9����fP�@n���Y��],�E�����P��Ւ˷��۶�S��M���H�,ڗ�m����E-�e����T�ܺ[V0iv��X���	����6�sM�f8UP�!*��YGvn��S�XI�\��e=��eLA�����wm�CnZ������욲Ή�#2�������N�ͺ5{ݧmk��N
�bXX��J���/J�#'�G���\1�n5�$�"��S��m�I��C�Uh�wr1Ss\��!/X�̫�N��e��i��zTce�oI�q�%��A�0䫔M���%lЃ�P�F��v�Y:f��Yt.�G�3`O͔MeE�#��^�-*[Q���!��Wr���ɵ�z��l-ef�Z7Q���h�b�AxN�o<6�����px���US�x�9��T@���E����y6R̤$�kU������W1�1���Ou�V���I�3Wn���s�C��k(ʦ�d-�­��l��0�����n�3v�����L�7eS�Okw
pꙚ�������՚a�2�{$��yT�̄����$m��#DN`�m��t!�`ڭ)˽O�y.�sn-�E��t\�����.b5��.���Y��[q54�/u��4��eDHKvK�>�bܺLǉ�u�E���5e0î�N��t3u�^(�@_4j�@aà횭�M^U�7���"s"��-�tQ�L�T,9��[{E�[�k'U���Q`�r�)�1<x�o%����-�;{&\���"�z����|�@����:p[�[�TUR���@�Ǡ�t�Ǯ�y{�+(��	���8�,��f�4�Wy'�2V����V��%В��e��#w�8�r��M��WB�ˎ�mBJ"���[�%Ս�50`��$�NPb�#q�ݗ6�j<9`����,w{J茭i��KjYY���r��ͰTwJ�^�S.j�K^�a��`�׻��n=���;i�xC����J�Y�CRq޹��.�SV�\nZwwUj��Ź�+�n!����k������ç���,R��e�$f�܁^��!.�v*�3�����Ǎ]��cmD�6^f��1;ZjU�ۇ6��=W��-�{����)�q��z�Vf:�1�yo\e4�Y�����R�ل)����&���ڴ`y���#d��e]:aL�i�X��L�4ϵ�������yj��^�IDm�Ij{���w���i��E�#2�[�{��P�Kul����ʸ�λrC��A�c �l���8�Sm^�V[���G/U���cF�Tg0��1B�Ƀ:3YW�1K
�z��t�WGd���k��Ƕ��u�S	�U���J��r��UBa:��0v�ޑ��T�=��VL0fݻ[�O2�m9����d[5{�ر%�[���ۡD]V뛁ŏ1F�5��M�e,R܍�JR�tލ�Hڧ
ASNf`�#kB�@b$�W�ȶ��i�n�fb��JU�Lɖ�ڼ����Wx�34�Aл�{�!V�7�8�^)�kMҺe��s�v[kV�����e���LӖ��.��lmI�HU<1	�'tf�Y�l˷m뻟`����N�5%C\ڳtk~�>a@K�4-O�N£����?jWoj���N�ط�����3% �
́���Te6���Wz���b-������bKj�Q���:w�d�0n�D��5��;'c#k�k7R�KC2���'Z�KB�˱CfiX�i��K�e1,]e��3nF˱z&ff;���)�.R�b1�Ք��{�F�Y,UU�U{3q�B� �$��S�WV,㷟�w3b[��Ok��{��\�x�C��wW��Y�u�l�vf���SO�h�Y�ۦ[F<Ԝ�*�M��%%*�
���Yr[�j�RZ4ҭ�S0nY�kR�P�1z�U�U
���+n�kǎ�يX�>f�O�T��Yì�Lb0��U)�X���V���
VIP\�c46uj��0Kٿh�/$��X�N��fViWXշ��Z�V� �i���{B�n	�u:�Ն�떅�NIJ,��rE��5�/��M�*Vi�n;�Ɣy�����B�p$����V��1P:��є��2��d���Ǐ+w؆ZT�Tx;���TvJy�FK�@bx��ô����ܥ�dĲS��u,���pԹ[���_-�7Y���B*j����,L����n��ǰHhd8`&0����gXy!ߥ�Й.��lY��xr:��ou��L�U�)�ݳWP�6w�d�m�n:eF�a�Y�C��)�.`��%�Q�t!@q���K��r�0�K/�?�q���o��ŴBo��Y���o.pjo&�AfR��2�YWR�U�U���!3sV�V,�\ڕ���flնE�(J�z�2�0�xǹ������Yͦ֨Z��U^��J��b��;CV�Ah]Rq
woMBm�
��z�ts1KpP�ҺYX��sU���eѻ�Y�Y��*�R���?���7����'v��_50L���u��6᳐���k*ݨ�B�P+Ue���KB���=ׁ�bVw��1�ʹ ��☃��.��V��m�֖p�<6^0�-�jL͵h Y��^�	6}N�=���x!���h�Ѝi�YD�,n�ZY�/hL��I�v�ָvj	� �)���F]HQoh=��Ʌ�Û!�՚��ť�Ri��щ��ʹ/-�;y�Bژ���hHc��nL�{�^��r�@#[j;a�7M��a�kD�zR��a�f��:Ƙ�KF#�3$�U�Qx.��"f�K����B����"Ǫh.���G-ێ�N�Rbf��7��V�*��{NhaR�@u�ǌ�̫+;���X�Y�)2�[���U��lMd6�[gmո�Ȉ�ԇƮ`T�m(�k&�gj��]��PY�V�h�)�� �q�˴(�D0��P�Y��fb�U4��dh��JZs^�-m�R����Z�Jёnd�a�	�K5z�}m��Ih�d]�T�jH^��tAyN���൲�^ő��I��*
�ӭ7zF����<H�ۭ�U�!ٚ$h����b�ʵr9�hB2]�a	hf)Zɨ���`M+U�a���n�Zp�ۦ�����;�n��:��3&,)cl�  ��7�ٲ|�H�^��jK�c˸Q�{�<��'֮i[��,�БcbD��#a�ɢ)��ͫGn�Q:�4R�I�x�ݵ(3z�R��`a
Ng���y ��1����v��������{��f���nRV�œ+����&�v1���X����W��*�nC�O6fnR����N&�܃\/6V	�V�Z)�E�R�7�P�.�t��Mi[������3qP�uA�b�ZFXea�p ��8�:H�mEd���1ۋFa�)�ٺ�#JV�ˠLٷ�)��h�*�9n��5���{��Ff�a��J�ѧ2�,l�/U-52	�`f�W�k�;;��,n�a�2�ҡ��[�ܭK��^��*EY"�Z�QE��G.٨.ju��K�.K��6��z�B�Q���Qj�eҡ1T��^��ŤQ��5%�pXBXLSE;�,!Y0��������Mr�T4��t�!]K(Td��\H+��#S2�*��i�&f87�AD�r��-�ZF�P���.��oM��1�{Uo(2tֻ��4dQ�-��qw"�w�cu�*����3C�fn�F��6�bU���u�\�ñYn���asM*�V�JE9�xC����@�ܓ,�0[� K��Y
`�fm�J8��+N5h'^�`K��+p��h��f=n��i�7�A��6�H	˸�l	[b�`�m����ji(�����yfG*�UD䯡̹c0I0���L;��6�b�+��8�w�����C���U����q�C�6B����U�_���.!��������q��9 Fg���
:.��)����:;�ԃq�T�������6��^WI�uU��\fwY����ׇ6̳�rp��-����{�(_�8Mx�8W.��Ia�6�lr��g:H^�އ�l{rT�d:�ۗ��=@	�wb��si۞����;����CF���5�Ue���1筠��^���G<��m��דmӃM�ݛ�W�mm�=ے����g�E�[<����v��*�v��=ZwW&ۮJȷ	���͍����<s^6��ݲOm������X+���X��a,��,KX���V̪q�W[5���c��8�y�	�N�p�6i�J;n��틛���#���/=�u����s�q][����nkkHU\M�3��v7n�����p�q�{6���-��@��l=�7��ػ:��hx��#�����/%�n�l�n4����I��Ƨr˷U�^2�ϷB�R[��l3R!k�۵nV���oG)B�Ͱ�T�n�Q��ц�̈p�����i3N��G(�1c[���L=�i�	��S�Y�[P �g*�/*p��Z�ܽ��>�۔6���]�x��:wh�[='e-T>�Ҍ�q.���X�vz�lY����}m͋c]vML��錷�5��H[��|�Ҽ�zB�%���v���y������>^�'���V�k�.���n:��m��/�:�ݸ���*�<j��/�.����u�'�y�H�v�kk��$��u2�eh7$�)��׎��yy�{c�K��<��v�����*P��7�,o8�m8׻m>[�ۍ{8s������%J�p���8{���<wn��"���':�u
�����qw��O1�;����G'f8g��)W]���mI8ǁ�ݮ��Lu�݃�8z�a�d�-ۇ8�����nv���v��F�:�n���,�V�;`k���Dm�u��M�Rll�i�O�K��^�ZA���v��g��b�Im������t����ɸ#!�xF"]U&��ݥV2��&���vt<n�c�9e�m�Yp	��y���Z6}�m���pĮs�3����u�m�'�tr:L�´��b��\���Of�c���ݰnkm2s3��6{q�v7iꛊt�nWR�^J���b���
>�F�ӝsm�vq���&�G���1C�=]�_b�U≎^��vx�c��='n�hP�a{�qcA�����ݍ��Ý�s�L�z�����d2bVc�]Ezے��>��po>."�7��6�R��.6����\ս��::c5�*;oZ�au��v�����n'�����5#fm���h7��8�蒾7}��ҚN"t���55�86��U�v��{�-�k��`s�n�v�� �ҹ���&�f�wm�t��3nMn;c���+��z:�z{7W���pq�f<v��cs���ۊ#�m�Źo\���(�Lx�k�)�����3���k�'����smc�n�+�ܛ��3<��L
x��n˺7n.���s���m��$ݺ��;���GEl��G
�z6�ٰ�bH4�+�wbN7�U��q�r�i'�m��#u�����:w�F���dF�9��k;��csj���6xNv�ۉ�Om#�����:�P�pRcc�qu�˚��[k�}�}��Znv����*Sc᜻���8M�x�%�/�g�s�gq5��.{t&��rq��C�U'���¡��aXv��[���Xݓ��جh�Ӓ5��s�+�!m=Smtȧ��{:s��y//p��kj�����۫�w��i!m�����%tH���#�x^^1p��Q�_`�l6�N�s�n��nj;<vu�,l���P�n�7+]6���[kwM�t���L��筋��4�mz����\q�k[��ۉ�n2\���)���ܛ6꽹s�����vv��^�1�붘Ɂ�n�����`�mڷh�\)v�N�vY�G듦�l��n�K���_v-��̢unzl�qnU��î��s��8�h2&ƻ�o�e㮋�۰V��9D�F�q��]\n)8ܺ�Z���
J���d�Ş�IC�Ηq\�P��-�9s�QOs��Q'<�"㴻�$���`��an9�-c�{\'g>�}��
mZ���Ș��׍��ӻQ��q�:6�'Ey���'[ۖ�:M�/g��ٻ��]e�p�ڤ⒎�eru����.՗s�΍h7n�������&��ɗ�g9�d�8��n��B�:<�N�]L=9�.�2p�x3�t9�omv.1�\Gmm�ڗ\��$t�\��G�Ol�k��m���w51�w��]��6Y�[Vw ��e���^F�hu����rIC�;o;%���DEWk�uomcN����4l"�o�=�8�/*�vs���!`܇�k۝c]S���T�c��$؍��\SI5�]�֒냞�
�c�������rv��Y��m��<�dq6yu͂ܽO�m���l�ON�.�V'�\Gd�ރ��4\n���w"��C"z��iFK��D8n��6+2ێ�8��h��'nق��wa�#srE=��#]r��cvq��'m�gDZ!��C�>������яg��S�q;�Lr��i��Cu���&XS]Z׀H��ݵ��-�Iw �v�$lgQ�'j�j�u�
��f�ԝ+����ۦ������[n����@��,��K�n1C��8u���`�Nغ|��w�b��a\��b�m�[H���;f;l���g��<�\�h8�zՊ�{�l9�p��vv���q�e�U�؋��v�uU�Yy����ehm�͞[��{)�G�a]���7e�n�y����G]�.dw;��9����ͺ5n�,哷#�.ay��3����9�t�v�(u��=h��|۴gmv��7��h�-��H��]��.��K�
�n�3k^����7`@�x��r=`�b���v��F�'�K�:��;`�n:9��n���&���2^B�3�/T��.zJ<�i���(c���i�Z�ۭ�a�4vl\����0�%��s�V�a�]1�2<���p�ϱ.^k�;�q�Y	�,]���(ۃ��㷁�5�CeM�b�w`��_-<ghX�!��v��۷Y�TD���..�ٯZv�u��7e�g7���ɳ���ŵ6���n܍W)��v4��[6���nwl�r�Ӯ.=<e����dw	M�͇�6a�kqUM��y;�	�u�������.Bd.�\�w\�M^Nh󚮒��v�ٳw����%wV�p�u���v3ζ���c���0���̀<�v�b5�ٍ�z�sK�����t�R^B�r�`ޞM۞��н7G9mr��M>�k�kKx�.G]\��s��z8�͓�G��Ǝku{[h��.G��皷[��,���Ts����^�6�۶���zlm�.x.nv�w]n�%t�Ľ^��B�']y�Qe��n����]�ڷfɮ��-�;����ḯ���w4~NM��˸����G�#�뮸�{�h�d��Y$�ƹ6�!�6�k�'�4�͎�.���-�����[Z#������8v����
㰭$oj�ę��O 4SmtOC�	;�wnm�ڈ*9�f��\�L�v��G.aݽ;p�nʝvŎ�lmPY�����|0��;[2]bK��n��1����X�>6�%�������q�kR���M�I[YY�ZR��`���>8x�ș�x�.�O7's��R��\����l��M����!�@&6��:�n��"r\�D�k&�8^h�8����n,<]���J�Zmȸ���v9��y�WX\�n�;���^<vG&�NXP���Z탗��YC�W;�6-���N5{ h����+,�in���ڍ���dx��]�x�����;���i�*���1����D�jCl-���>��e�J\���T��D4�WAsیygֶ�ݶ�u��A�{a,k�ַH�3�V]\�-�61&����h=��0��E��q5=\\'\�s�����nz�m�\]���q�3Jv�q�ɮƚ������g�'k�YOv3뫎�
<IA��d��s�ۄ��7b�695�Vz�h�$�k��e�ӗ���{Y�[��C�k��w$�]�����͏�x�5=��n؅��ݩ��޸1�Ş����]�q��8{#���e��n��=ڍ�凱'���.���^�vNV��֏vWe�q��mW]��턳��)��v\���7f��kB��dA��<����v垌]�&�';G$����n�mθ�}p��ю��q����{y�kko[�׊ҽ��6��t�슕�z���"���=��=�7U������v���|��ݸ;�^�<6zp�u��,�-OC��r��C������v�@n��-ɗW���L�8c��<�l��9�t�p�k���li�v�pp1���h�6m�G����n���z�^�J����ζ[����;D�]�ͫ�keJt��v��A�����v^�������l���Z����Χz�	�A��v����]�*v=��=�oK���#�if�4[;`۷
��\vcq��7����{tF�5��H܀���Nڻ��Nn�7Olv�g��nV�G&�~g��m����|�Wm�anܳ��9�����ŋlc���s��X�o8�l����S�0�E747<k��7i��7c�I.�<+�\���Rpr�[�L
]��fv��=<;	ۭ;��:4�On���WF�=�W������\h}��N>6�lskq�k��1k���/s���Ѩ99���h�[�[�w�ǎN�(v�I�-����G%�ۇ�-�����8�䶫�]z�;��Fѣ#�c��Fz��`5���mDrp��֍s���v�̙Q�z\۝�p��=ng��brV^v<������빿��?�f fa]��pi���g))T�/.�V�G�q���ٶm�>�p��a�v�rtm���X�(�EW�R�3�ٺkXI�v.��X���s�vĥ�5tc�do&f����t��.c,�h�۟�1V{��I�ߥNoO՜�7����=r�t�Һ\��^�}�K]���s���~_? ީ����͕SI���4�g�p�p~����q۷�<��3������xM�qo8cD>�k��l��stN9B[��@�*�Y)%nM��KSx4KDu���t$6��fVsv�)FH�*]�BsH�T�\���Y�S���-�%�IoR�^*CSRɠ�T�,��5H�6D6��08�nG��8:F;������&��O��@|�{�|�N����/&����̂A\�֚^N�]�-�V�J�R�7Fd��ߛ�Y:���*~�?f6��cs喡J�&�(���%�a͉���r�n�c%��B��/n�9R�u�!�[~nn�r��<u�=����ó��|���㏎����D��ӻ�mt���l+"2�9�7g��	d�������6/`������qt(��_�/&q�D�ZZ�����se�GE�/vܓe��߼|o�ȇ��<`��#��G߅���9�<�V���Mꢨ��	��SF/�s�K��$�8�ؕ,���Gd��;�(��Q�^����9����E����f�'RV):��{��9v�$�l"�(̊��u���͸�>��|v����v ��;�>~:�e8��M�\z�J��*��V����4s�^�F��kȤV%�I�}�6I��D
&8�D�uN:��ا]��TynsI9%fH^m�'.���\=K:탍���wߕ���e�$V����ND�I�y7�!d��+ο[��q�?q�p;e�Ԇ�a�o�����be�\��P6��-��מݕ�wڴ~�F/gm���vá��-���-,{����;�r�����c�m���=.�wv������X����s������Z=kA�~�K��>/�6۝�{.�ߏ^c'>�ɐ�o}<j�T��� ��	�Ԛ'%��z�96ݥ:��0�^m�awί:�)Ya��T�Pt%Qb�4!6���;jW7�)�
tn�v�Q��Y0m����ѐ]�[�����v��R��ITf�FW���]��P���M�r��~�N�e�y��;ܡO.Jr�R�I��#Ò79f�lN۳f=6����Aڑ2�顸�W��H��c±%^i�iy.R�+
\��9n���uF�r����o=�nK>�D��-�Dd-,����NyC"񆗳=x�>N�;������r|չ{�#؎vM�����^I6���8HRB�mʯ���<�;��*�17�4�m����6B�5wK�[;���a�)ۭ�O��>��Y�����n^N�=3g�aa�7�Q�뜐��N�h܎28�AKpc,fˍ��{���J��=�6�*YcډUAd��s�e͆���H�!]��U/n�q���*���9&FX�m����s]A�R6�I�%�q�Yty7��vګ�Y��񯜟/�s���ix{kuq������]�b.��Ș<�n9y��e��Y�}��c|��؛o��b��ǆ�N:[MT�.�,�ˋ�$Hڮ�)�c��&��7����}	m�z���%NТ�������dB�/%6)��뭼r'$*'W%�,rR��[�d����j�)��m׶��Y#�F������U�Z��݈�$�K�*�,�9_���Xp�"x�n0��nkm��P�(��Yw�b�V�ͼx^g+[v�1H���9�ד���Ɩ�G�U�#�1瓝ʹ������QT�$"���(9�� ����4l�X�Hk"�!Fތt���s�=���\c�T��E�f��%e�F8�%�ucVK!c6Ԣ�"gR�rL�j��>6�Bf�l�c�ٶݟn�72ý�o~n���;�f�NXKF�$H�"�.�m{�+��^;�������ޣ�Un=���''I������|=��n��n$�jm�4Mu��kZ^�c�p��;��5Ѫ��ކ�a$!ܷ�5ݽ��s�����#��0�X4�\D�2&�����n��=�cy��|` ���K�ۀw<�v����k��&��L���R����˵�QVq޷BK���h-z��+k�&���R�7v��Co�MC�u��GX]���hѤU��Y2�%��\ن�Z�p>�qD���n����^���%X͉Ԏ��"賤n;�#�Fٓ��]���賵���VYN]�bI��KR��e^3���wζ'!̄ͷ���zD��e�Y\�w�l9Yޓ���:Hs���T᳐��sEy�����,���aPP٬˃fҷX�Q���im�&Ɋ� �jEl#
.̔�����{ܻ������R�m!Fl.�be��7E����\�JBI+sf�ݾ'����si�	���0f����Cv&��4c������v�3`਺�ܵ��Ȯ+&�l9Ͱ�)'l�W���D�r�[-c;��
G�jTF̤ۯO)���͢�I�X��&��cۿ>w�_0rm��c����ݴx701�����>�tx��<<�����o^�q��:��o�.��6(m���tI5��H䭬�6F��6�=����m�o�1�o&�H�r�T�A�ki19d��h�n�gS��W�l�E���]mNC�W���'$T���2��F�kuhL��{l��T�azz�8kal��,��'�9�/wu�kX�H�ͱ�ȗ��u���7c�>DQMߓ�ۋ�%b�!Y'6n��sf���\�H���ܘ��.��ϐ����n�$D���2�wpR�[���Vt�&�,��LZ�ֹ9"E��x��ַ/;��,�a�%ۭG#7��"ubηz�e�v�b�C�y��b�ɻK�u��I]���Ǔ���H�Z�e�4G�-H7Vv2ږ�ń���##I-����9͍V�޹$�il��9`렕$��+#�!�0�o)�W^1��h���KcM��2ѥE(�3��s�x�w���=�wZ>�g���݋�;�����v�:�˜HkW�᱑��-�I:H��
�
�ns���>x{>k�B�F1d��R��&!X4Kr*��rD������Q�T��*�!.�{�u��ʄ���Mb���n�~�����rt,z�<��N=n��Ŗ��l�&l��$W�'"$�	������������_��"A�%,���!�,�N!���k[�ck#��˩Ʊddd�����;���@T�{���nm��I,朤n�KqK\C�7�9���\��k�~�d݆�z�]�-ө]$�ծ���SK+q�ݵ�<xِ�^���;T�_n�ٚ�\��UG �m��N?z�[�S��ȣ����EY���7��a:�j���y�{�<���G|9xȜ��x������kUE��܀�ӷ�sc��3��j2��^2�bT�l�E������mrŤ�i5c��]ay�w"�n3d���V����l� �6QDњ̶ƣdR�"8,������me%�[��JY[`�,M�;lb0��`n��-���$FB�Z�cԇ'8M��\)��nۤl98�4�ɼ;n;G��s���>���V��r���*F*2E�F��Q�\�:�R�X�K�K(ճ\Z�o3H歑�#Iq���RB[pa)H�6@�����[$�rK�57HA
)A�I!5�B�M���5�ܕ��q�Xw-����vY)��Ȳ��Nj�,[$cN0��`�ێ�4�9w�%����ƴV8�m�y�Q}�y{pra\m� �pol��V^nmIB���l�ՌYMM6@`4r8DLҒ6�ʍI-��Rue8�(��$��r%�8o+e´�*�Q��:�Ged;m��>�y�����>��s���t�wZ�냎�E��6�����2��t��J�'#!�^]���,l���e.YHR#�c�I�D�dfM�Ȃ̓��Mfy����X�����N��N���"���,��9#�q"�#)msZX�b�R� ٛ,��|�N��T�d�@�����i�7�k�D�ͥ�⤎δ�Q:���e�i��ّ!lI!	umԦ�v�1"�7ae��,Ֆȣ��Dd�A7f9_9�:�7m��f����s����N7v)�5��W͔�"�rNl[%V%�]q����4��7���X\aW�&��$#���zz*K%����Am�"�גh�ɜ��Ŭqg9n͐`�+�М������۷��嗢m�c`��qcm�o�?
��ɾ�8���X�d��&YcQ[fY����V��ʡY͙k�u�C��K,���\�Ŷ�I�ٝ&�MT�����wn�-���ۄ��V;�"rJ�h۳El��r=�!݇��؇.��;o�&8�
D��[b(�eE��;>5�c���n���/n�2��S��m�}�q�<�l�U��t�V�G"���f%���I'Ziv0��z��jUI�\�����,j�c{RN1��*IKe�l�jҥfVDd��kiSR.�X���m�:k���!�M����k�+1*�)d7b�HJZ*��F�E�ٯ65c%�{���L�;�{v4U�Ƥ��,�d&��J�9�^�r카p�KdhH0Y�˔�$6�nw%�9	 �A��*�9X�E�8�ͯl��dVIK�Pc�aY�V�f$֔�*A��ZJ�ZԶ�G-��y��
KԂ�v]I��AE*���
��:n�۲e�Y֜�x�ZVU�m��d!"�6���:>��~!����c�n���㴗D�K"�T����6��AJ:�!l��Er�l&ɲLc[�\�G���Im�9�T]9cR��֜�b�Ke��DI1�2�����u5�M$E���b�s��i7jf���I�Dm�\�ik����Viu#�+�;\'v���D�Bf�k��4E����f9�F����˺Y[���0Ԇ��dr@^���d���y;|�^w` ��s���f�<��}�O<q�
gt;gݾ�����xr�[JČ�݄�Y1�]�*�a]jk�!E�6��ib�[�<n�Ҽ�#� �J���L��;YCm�x��y]�����~�r v�������Ib�1�Z.Y����"����4�Dbd�K�۪AR�I$��*���;�4qr�ɖEm�$�E�N1�A��ʱ�(ֶE�_%v@��:���"��%��K��I�H.q�3Q��rI��n���)��k5*�Ȱ�c��;`�ce��rb�
HU��Yj�`��W,�d��$Čdb�HZH�j��Id*�h�1/|t��=�L�O���N{w8�6q��0?�a��a��8����32�`|n.+C�1���vO��2�kU=���wh�b켓u[\���ۭ�.`q��Y�j�<���#�]�ǵ�#�GUmv�n֭���s�m���V�Mi���8,.��R��i�kss�"�,����J^�m��.�����E�/F!�F�v��Wg�����뛨�7�^;$ԝ���a��k��jv�����#�y'��.�\:�,��m�d��M����k��[� ��d��&�Ģ�;u����ζ�ѽ۱��z���!�n�zؖ�M��7��v�����+=ZB9���t�s/��U���Y�e��ٲ���ۗ�y��`���OE���s[��!ȏE���`��Ƃ�gm��:�u��w��-�z�:lmV��լsA��fr� zP��7�����@(�7G�� ��"m�f��h�v���#:շ<�09^y5"��e��aX����i�5�.<�m��5�\����L���5�ݶ�k��t�W.``��Kv��.�'κ�p=��a,�F�	mRہa�vێ�ͯO�n����֝���i�\�N�4E,i$���a���F68;:����C�!B�+�3�ny6�������gj݊us�=\2]��u:�u�Ky�	�=��1q�۵�ݲt�5���^�ع�΢���t�y����u�E��n�*���z)�9����ۮ�� �\�1ͻ[GjYWI��LK;�r�Hm�1�Su��e���W��Ȥ[����`��Tܻv�G��r��r/5�����Ԗ�t]��n6]�z!pn72��n�zT+���q����A��]�n�q;nޗi�"��q�/;�o�����&�(�n��lB�F�x���a�ggT�=&J�"�ˁ������m��������;o���rOu�Z��bM��M�J�&���v,-�<���q� �W���z���p�ݶ�qt��;�97�k�[�ے���d�Yn�k����i6;����9�	yή�lt���u����y�\��\	����d�뎺������L#�'n�;'V����xv2Z���gz'���OZq�;���3�KA�m��c<�u��:�C*�ۥsf���)��Χ�vz���tg�ˁ������5kr��;[��ۋv�XR�6�v�{v����EC�clh{O�W�:����zew�����q�E�d��h�,Hˑ���,(�!��e��YiHH#�__%�������p��/=��r/"U���@h�[�$�;:]l?f�sW�W��R�]⁐&R��˂+^�ϫsa�H��kn�2Bbm��%�-B��������qfz�{���Ô�_Z�&�D���Q0I|�jخJY��3��� te��X7U�]T)6�V�G�
��ZA��qfr�]�+Pu{��Q"�H�G
��(a�5��,ɾ���c�rVRw��� �0 7���QC���J,����DȊ�YxoCxWO,�2��ƀ�o=Bh4Ƭ����Fs|vq��E ~����*�Tj@��ir���!����tRh@�e%����?�`�\��i��Ʉ��n��βU�&/�Θ�#F�%��G���#oNd4��R2�>�9|IVu��	H���p&S|Z�^�f㣰�qb�T�v;p��'i�Og�\�p�T�!G��d |7͟q�zO�?tߍPM�w���.�"���Y��eCLG!���D�x�^KM5�=־p�Cpp!���0��ݏ%'��{��q��f��[�����a"�q�vf;�735CX�s^.��M'��K���խά�{wrUaQ�J�ފ}�^�WU�;)v]Q�=_;�S"R��l���
�k*io���Tw��z��lt@�o`�B�n�49���`%���#$�W��t�A��V���n��M�	����;��j/�V��u�� ���/R�ZL���z��?
ɉQ�PE�#��L/�;�g}#*&����2K��:�,�<<�ɂ����n��(�6��$�vj���'�G���~��##& �)����#^�"�l�ԜQ	 ��xTD�����^��>'�$GK�djD��]����u�#�jhn�S�_a<m���3����Z��Q��@���$�E�s����BP����q#$y�P*�=���k�Hi�#��[�Cr��n-[=
 ���4n�ŔY^��+�f;�3mن$n��7x�jn��l�d��P�u�U袙ϭj�έ�jƴQ����hq�Y#ǃ�-*.Nr��C6��0V����@!=����Ȁ���
}�j��.����\f]{E�ͬ���� ���'���;�#a�	p�����v�QH�8��
�S��1<4�]�ח��B�
ǫOq*�q�Q�zKP�CD����{+D_�����m�)S�XJ�Wm�a��������ѵ�}՝{��mi����c6�7^�^n�8�e��`�}�>K�n�����o��1��`� ����U����Yk7΀�.�-x2(��@ګ�z�A3pbzP�R�{�/yeH(���j{�IA���@�4�Xlh���G,HSN9*�+9W���͵�_ù�Ҵ�<�CZ��M���C�
�ʴ�)�p�c��郞��m9����9��	���ݭ|A����e4Fm\���ŕ0���j��Y��v�ٴBu�<m���i��u��k��T�!���a᪢#/�3�i���Ӻ��L �]fN�:aB.�f�^U�+:z�ڸʋ���_�,"�ZqD�!)�v)�5�g���Z�Jk��+r`�+m�E�����۱9L� )�6O�{����`�����P��%���m�e2Z���V��&��[Q���CE7S�!�묯{z-�����F��wq�CDļI�!��	�mh�� a�q
N*��N5t�Y�����b~%�!�2B4l�6{�]��,$.p�D4hĩ�ֺs�ܾ�ݭw#t��r��T�q��i*�:�{)��e���Ke��·���'^��h'�)Y#D��f�S�7d��{�i}�*�-�aZӟ/����X�����-(���䬴4~���\3���N��1��##�}͚g��e@�	�Y�P��ծ���!����;�J���@��Z��8��E{&u�K��]p�˰gN�iU�Ex�{[(e���br�֛t�*�߅="���~�ʕ���#f�j���0"���qM��/5������<�eX'��cƈ~������I���z�d�2�Su��_/�{e��h�=[�+�e2G��r��v��=%ـժ��#���<M%	�a��L�'�X�Ӿ�P{m��\2��9{<΄7y��`Χ�W_N�J�8x��l���N��y��?
F]�kkX������&G"�s��᪬(���I5ݢ�F���cAxTV*p]�EE�O&�YB��۪»�;I}g�b:�$3��O@�e�ȌD��`�#��^��ڳoϦ1����Iz����>�*�����P�3�͓9<P
]��8�#��ȀqpS�7�Os�L�f�zl�p�KW�+�wS[�E��~{�j]|+���z��@R�}�,�zv�e+VPv{�:t}��\�cn���������#iAn}[��Ѷ��u��؍���q����\�|&{x�;��\m��ݺ�Z
�N�N�(��\۶���G�P�=������㘳v-�i��Y���:.�Z��8���;��,n:\'�۟N�#�M�lƹݮ`��c�"�c�t��0{g��sp��Xg)�v��f�u�v� ,�=u���G�\C�)�����7g�vmYqu�66����c�U��w�Ѭ�R�`��?c��R�����γ HΥ_���ӒD�L�溮������O?W�#�d1�z���Y�NVdU:��<�l��t-#�H+�!�2\i�[�m�;��$4��W���T.����gK�9f�H�ĠR��Nj�<V��^.A�C��˾��دO��Ӭ�t�,�<̽|�,%��vT�O%��/}9!8ff��~�4�y�Te���;��baU[�)_=HFjٍ
�q�$�[|V��>E�[+���[pe��l��Μ���L`yQQ1���SLdӻ�f���`��P��rR�D,Lj,��%T���0���5惤�ӂƂ�2c�0�)�>�Q}XW6�fgt�zt�Yi4�\b�[��q̷���5���Y��l��$�Z�K���i z�`�]��E�x`���M��s�#PY���YY���s�S�WK�N�q��Zʓ�j��5�a�:k��c�̙��:�k�|:��,�SwAf���ՖQ}�-��6���8�U¾�r�\K%v�	!"��Y,gg"Cv�P��l��OJ��#��J#�p���;�Zr�d�#������]�u����l5���n��+S��ˍC[���z�w��AI�fzEM�tTɰA�)�N�i�i7[��fz	q���(p�։%��[��O���u�/%��u�M�m���Ŏ�E���B(��Z����鍊�t%Vk���+⢑4V�|��d9|�G6�Ӳu;�«��L/Ӕ��a@��]��<'R_�ݐDN2ˈ��p+��ξ,c�湪x4)��]�Z����,7p:�|��Y���L�����:��8y���.�~Ē^~�2S>��('$�����)�Sӂ�>$�GdLW\�WE嬇����ᣕ�W]����
O�2��b{�Ξ�h�KR"����v�g�4		��M�$&)%'u�Qv�n;����A��s��%�F6�q��v�:�d�FGB �H�D���]F.��`�#��Ad�u�R|���}ێ�l=�VHd�!���*��zĥ��N�:�ҽ�r�TD�	%�V,W\þ_�M���.����Y�Qf��`�:�U�<Wą�'�I��b���*s&
� ��z���]A���3��H�\�.I,�8ǎ���{W��8V�,>��-�ץ���gZLk��Sm#%�㚹e����pX!N7�J��՘Ru(�|pmn [�%���%̉ͼp_Sוp��H�c�V��	�M�b+=]eeC�ծ�}�+���$�{����~� �D��R��$��$�BL*E��~'Ç{������u9nP'h�I(��->�]����,e��9�x^�XX�
�ؚjb�S��Wu����Gp�d
"��pyL$Ӂ�L_ڭ�$�?�>��u�D��/@�Q~<�4%q8�c�,i�K�V:���:�C�jVψd_���u���S؝_[��eG��X�LQ�ӎ˭���eN���,;�̙�Iݭ͙�g^���Kv*��w󞺡qY���X�k�|cY�Og�a������9�6�9(!9u�����Ň�J�7�ߨ��H0�AEa��w�Dj�Y��Ꮢ�[IJ��V�q��A�5Yg�N�+���%�ґ�k��n%�H�
�GF�>��	-�	B"8�ǒ�H�ע�J��g�')(����vr+��S��~�p��k�j����j�f�h�i�)�e!P�. ㄍ���*R���A�"��z��"K��',�t
�F5{@8�w=� ���d���Ճ��gX�lC���f�*+��}R.U��n��u��f#7�J��A�][OK͑�(U���hfN�.�s�:rzN#��1���NU[z��}���52Z�aV��p?d20ԂAR
��I8��]�N�J�v���ԥ���ܶ��٣J�#C�K�xg��ǉ���=w�E�����ǅ�S�yZ�d�:+c�`w���rf��eM
�7EϿ�ﵾ5�j�fn�5ْ��X�O��T�c=����W\@�1����(��x�l��̓�^�ָ�c5ȫ�<7Dz���R��0�÷O��nB�rT��㒳�s�!����oh��e����<<,D(�qn�o�B�UE�$�̃��,��5��b���|`����8R�a���hW�)���$"B6e��l�C���VA��3C�#A^���5��%�u+:�~�����T�����1��/9���OÒ6+N�$o�����q�e���dh����'<k)eУ��r����5�,�f2w����b㺦,����Xf22�4�s����v40���O����Q¬Z��5�Ӳ]�XX=͜]\��s5J�h��ɴ.7�K�Q�I��ys��]eȌ9����x�l�}Jtہ೧s�]8��`n��Z�+�����GJ���)���*�C)�
����dDT�!����]��\Ŗ�{ܿ���ջ(�K��]�8�{&N���5�c�_�Mʯ�8�ͮN��']n{yfg�us�6E=��\�a6=� ����dq�5�8�h�W=2�v������n[s�^ˇ�t8�}���t�OYy���b�!h����7l�6�M1�ނ�n,�y��V��<�s���WI�@|Y��vp�6]����l���z�m�-�����q��Zqv��c�ۧ+Ȱ�ncCw.H[�@N�����_i����5G�zU�kS��cmD P0��i9�/�zDۦ�~Xh�΃V�~�+�7�C]h���E$�%9�o �ì��sd��U�ƕ'�4�.'z�����R�OV^��0a�:��6Vn5yWvm^
/e��Z�bFD29+[� S9�𑃠`�f���I�ve^�7�]�Az�v��	E�sw�P@�l���7=5h���/��F�\��.GG<��׭�9�6õz�-�0�dР�U�ޘU:"x͞E�;��J���4N.2�K/N�={a�l��Tp4�d"\M�a�J$rǎj^�3���T�|�,k�z#Ƽ�&���_AG9�����]mz��H|��Z<G���A]9�8��o0s<X8Ɩ�6����t�V��fgZ�+4ʠY6��Ђڭ/��A�zw&�H%��5��3� A��f�>\�>�y+r�v\�L��w���uU��6w���#�>,�aa�2�w�S��8����ʘF�gW����E�֥w��b��	�����VYn%]v6�9�uQ�������KwW1�!]u,��Ѷ��t�)�ռ�:"�-��1�p��=7�d���)(lV.�{{� �@5g\��b��6�9��3RN!��I
M c�bZ�ۣ�CR��ߕ��#g@X�~4/Q-
�ŏQ����ʙ����V�uWP2BD�s�/�|H2(�H�#��E�Dz������V<�o�6�
��?G�0�m���֌#ʈ/�T��Wn���M�v6#�C��ye`�1ʟVҀʘ��B$Ya"T����>��^��^����0�]<�Xҟ���]lW���U�L����@�!�U��,E.}�Ṅ	^� ��Hj�f8f��l"�k8�r�v�f;�����@`q������uŰ� �S�A ��&0�!�6���+�y�����3��u�Qq�  �F�H�AS�|l���na!P6+�-�瓌�žX|p����D�E�>��0ё�yw����^��l��n���m�&	�%K1-�r۴�<X$������E�U`���~=��~y���44PD�r]�M�t����Y����X��o(ެ�_G��>�#��>�t;�w��_�	�9����tiR?o]��1I��!x�q��N��Z
P݁jU����K�X�
Z��Y�q��[�ӛ�����{�~�׵��y��a֚��w;�I�����Q[��\����B�I���<�*,�[��)f1��:�lE���4�a�v�i+�h���M��m�ܲm�ʺ�V�t��t3
�D��<�k��u�en��ˣ[C0_mA�@�QY�:�ͻ�yY1J�B�R�v'4q��,��
�L9R��$��y�t�� �w�]����Wp���٦J�ʝ�:��D�O-ױn�c���X�ע���L�F�͎PgJk�9:Ø[ZPU�s)�_+��']�J�MSsD�e�i�n�c(��TqL}}Ր���ü doAX7���r�<	�L4�el-�6��Z���{��D�gKG��v��>V�gZ<+�
���������)	��Z��B	#^�*�U�;�ʓ�C4ˌ6��p��=�{2�/]���}��L�Iй3e�t��������Gc�u����v�9T�
+�P$h0'tu��g[;��pgN�ҍ���aEq��9���F^�1Xc��"���w1�4vF.V�.]�+r�҂��R&��f�ղ�X�Z����K�fl��Y�D�6!�j՝�	�H����u�(�yX�����	Z�f�j��Y*i���̖Q�s�X��Tޫ����[�L��
��=�Q���� �Z�ҷ�w(��J'LK�w��l��3�Ķ`{�]���5��|~���Ή�a�w!�"k���G��{xt�bw���L=���R��?9Q�3�<������p>�X��o�9�GL��J�u����x�t��ݛ�0��#��9�^��ϻ�ϓ���߿�v��c!�V%H����qAc��erw��]�a�bgޓ5��
�%OS*W�����������=~ٙ\�#~��ޏ���t�o]M����_����e�}�2�C�+�ນ\�x��y��C�g�|�ߣ��Y��n�Ӈ�>�`�\���}���֧�W
���{���3�#Ӂ�"g�#�nG�p�N7η�ӿ3'w����>ɕ;p�{p�����J�s:}J�~�}�^�DȄs�R���!�>s\�k��ô5����W�9�!�+��'9��0�&��~
?
]���P��?b�u�+^0[+�]�i6{<]l<��MT��;x�Wt�ZD;&B��M�0�]��q�������9�"ju�3S����T�y>��t�v�fx�G\��ބ^��\�X��y��aԄ�\�&z�#�QQ���߲���o�h_����#�3�Ğ�2 �n�U����p�{�=z:I6ֈ)��5�2u.����ɇ�̻��w~�j�E�v��v�ۇ���p�
t�h��nT*g���u�:H��>��{�����#��:E�k���;p���|p��z����_i��0;c�~�k�C����8��Ӷ����ɓa�
�%k��s����t�o�+�����G��?|�]����p�Z~Azs����S��S�]�Kd����OS��f
Q��|�H�QzٜL���>����G�'�3_\�N&����u��z����8x�s;r&!���w����?�|	�iր$�㿷�oY�P�{p�g�O\P�p\\��N�?_:�^}��p�3�9f8GS>r������D�u�_���7#�g@vཡ�:n��@�����>�۳�s��?8�S�:��]ç3�!��wa��K�sO��๟�߿o3�\?X`�T]�L*q5ǩ�a�Ϲ���
�����epR֯�}�����{�F�y�Μ�MJÚ&ƳY��������2;��VA�V��.��]��i���.���w����O{�����O~��8x�ܘ~p�gND�Z��MsS��=��������|L}�P=�y��C��L�\�*�g��>y��~p���?'�5#\���̎g�DC�������z~���8�@�5<p��
�}����gH.s���eOv Oߺ�a�ہ�&D��%�뿿tn��7�����MmU��	3�q\=D��6�n8��q���Tz�ڭ�r��p���n��~AN9\��p�?~��ʙ�;����3�R'h{ה8�/H|�9�k�Օ�'^}��v��D��j�z�J���!�1bz�l��	���]`�'߾?zwt��L=����o�aՃ�u�������?"����È�:���:T_��\ψu~��n[�ݻv^�D�I�HV����jaܘk�������p��_�-�:䍎}a�B"2���j��9�z����9Ӹq����)�Xb�"~@���`k���}�<{bp�g��2�A#��a�k�9�ȹ��
����!�#���y��c�|g�LL���3vT�\�^�}��?h黻�]֖�����?=��rrC;LԮ��Z}��9�s�<W+��������p��\�~��ߧ3�o[��X`�����'_����e~u�8���u�=��+�K��j(t�������O:�ݜC����u�|�eN��!�����p�Y�>�j�����y�s;O�p�X�Hdi��F�`aG�����|+�#�g~Lʘ.[��\#�ۑ<@���M�|�I|�O�:N����9�T\6�CQr��y���9�s:sښ`�r@@~���C�;�28�He���=^���>��,���1�C�HC���Q�3�����_��itd�����3�?Y��.k�+���+��ș�s��*L��+�p����ӜL=�~;�w�����<xI��t�B'�}�*dsz���Nt�����8���~s\�gv�jeO��ʐMO��3��y׻�v���,0S�|�{��o�t�#᠂)�HzQ=9���T~����4Z�b�ͽ]\��:J����9����He+ۢsO1�]�u�Doc�PG�F߭x��m{7[���D���"���.;N���6��nD6gH�<)L���sţ�2��C����[�m�Q�Wc�ہ�۳���o(����S۳�~9�(¹6V0�Su"nk].��M����I����+x��nԧcz�+Ƿn,y��X�|�,:u�=�[�>'d ������p�G1v�:1���m��ɜ{Y��% t��q��7A�,�b�ۗ���B\��[�r��d��s�=��`�%"l4V�]��uv笖Ӻ�D��r�B]�|a����1?��3�p���T����N9��3�"�BX`�n5�t�O7��/N/��s;��P�j(D�`q&0A��5���R�/�G���w��N?'hG\"y�dj;��?{�׾��D�)\#SP��u\;��O���/��n��$d�8N�Φ9�q��N�1p�>�>�_��}X��|�zf8y}�*��>qC����5*cf�g�s�NgI��`V8��n���9\��Nu��x`���N�.k��ȘY<p��#�}1DP�4}GբO��{E�����ra�L*z�W����F��7CH��;:�g�#�>��þ�$C��W��P�O���w��0�'��V'H��W
���~��0S<E#�VaW�d�[�=��^��ٜ���;�����u��;���r$s;r��<�'�p�z��.��:������7�`�ɝ|C\"D���վ1�!a($m�%�G��_2�oO������@���O�}�}��̏�@��T<0S������_S�8�ng�0S�"y��y�:C�Ͽ��+ә�ȇ�o������ןw�t���o�N`�������5�,c B>�U�������^�p�̾�:�p���C#��0]���"����3�T;L���V�m�-��.ټ0S���v�����x�gLrɁ�.�}�~8n�;p���hy!DI #�D^L����~�O�{����+�gs���g�<�`�|�\��P�2�;{b�S��iە���	�����w�i�2�@�OD�G#�J�q��9�&.|�VxS��c~Y��aH�Be���`Ѹ��;1��Ĵ��Y���#��/,�3�p3��5���wxn|��*sهoIĈ�0S�Q+�N���3�"�@;H�L�8ifg�w�������f����Nܨ^�p\3�R�� ��� �.��>d~��R�"?rz�Z��k�O?~wrrT�*y�����|���a�}#���r¢����J��M�
I+�8�z�p�ه{���ĳ�C�����}���G�럆믮� QC)���.:�~t�ћ��f�J0�DF4�N��m� �
1 U&�����Z��y��j^��?�|�F9����&gNT������ �"o�pP�=&~r��g�T�'��}� ����+��S�����
�}�^$?}E���Ɇ�E����@��p��������;��C�9��<B��~|I�E�f�֫.Ύ�ܮg�f~�njW3��(�����3�$�{?P���>p�S����Mp�W��T��8�N/����DL�~�pP��9P���}����/vx(��'�kz��|��/ٚ���f�*g�S�L���}��y�=� ���`�����8��t���s��s���ǨO�؝j2h��f�`�������	����G홫��-a�����7�<�8���/~>�k���t� t�=@��z�X.%=������� q>1
�|��߷���\=�<L���p\8?e�{��n{�<E�>8�uy���$<L��u��ɛ��0�,K���~���IsM�l�|�?1�J�{H�a�|�C\��l�������(�nW�s;�����@@�C.K�Ή�w�y]t��>��(��L5������W��)��r}���y���dk���$��r�ӟ�)��ߜ�?�z�\"go�Té\��O_G=uï��<m��������R�Y秔K6����
�vǝʝ�9Q7J�l@+��j�n�aJz�^��ܮ�ý�H@�2�q�!��O�y9��I���h��������a����p�O;���÷*Vy��LJ� 0��,�j%~8z��������~pP����3�=��ʘ/�}׽�8ɮ'�+��9�?^S>L��8.�οt_�N�l�k�tۻz�����̨z�>N�]s=jT�ZL��� ��B&=���`Da�P����9�H��Y��aS�߿hv�I��[�Nesl��0*�v��W��x���ȘY	�SB��".x�ξ�ﷇ�oܘ�3Qc�}���S��|s8�$�p��Tʇ�&�{dZ
pT�ww���n���~�H�}J���5���*S��y�ᝧn������ƿ�g�b`�K��aә�3�:��Ow����	���D/`Y���lr�����I=C�x�F�m�~2��t��lL�E7�̍	�_!:��d�c��L9C�vj����P�����>s�<�E
��55 ��w��o3���@��a\?8D7�|5�L<����1O���	�6¡���s�E˳X�_��~=յ������|�E*x�۔G����;�>27��� h�>�>���}�<��|�y��w!��.�N�q���u��v�G��O�}���/����k߾Ӊ��tN��E��G�ai���(��탋}�A:�����zp�Ar!�L�r�z��p����p󗯤��E�������v�3�ʝ86�"~O=���H�}��w9�9��g�3����G�x����9���z �w�P�<@$-��[0\���\<���6`�u�t�u	&8[E��6}&�¹X�=u�w:�s�>r�{�l���÷	�3��w���׋Ͽ_����?���<�f�L�8ui}��#Jt�G@\ꇚ=p�}��Vn���?<O���*9�*v�q�
u�*k��Tʄ��7�H=CyC�8G3^Ҧ�y0�|��<�;p\#��*b���V�����}��N=L����S�ߝ�x9��C�
v���W̞�믯Y���~�=s#���\>N����:p��I���@����)H˫�>Oɛ��p\�t�~�ȼL\�ʟ�?O�w��xN���{���Jٮ�v�W"&>Z2'�������<c�I��*a��)�p��
�����}9���,���<s�
�&
ũS �����t�g{��W>�D翹���㇨�����H`�^��6m��J6�8�ۚ��G2�f�P*x�>����~g�@�B,�{`�~���B z���u0\68�y痙�؁����� H���t6�봊�?��G�1�N'H��{w�>C�+����|�u3���/!����;����Ϩ���MB&?Z��+��8>����;]��#7g0\��G�dȍG�K[H��V׺�|Dx@>�"4g�w�o3��}�\����pP���,���߾7�
o�
�i�F�B��k�_,�O|�����&����u�TD�l(�w�߽������� ���5F*�I�+���Ql1�A���%��WlɓE��)�!|Fl�N��>�#��F(	*b��Y-Z�m翳<OϚ�Gο~y�{<sP�+�s��a����眢�.g�ܝ#��.�+�7woY�a�@�2'-�z�V�G�*T���/�?$��w�?'����ꓐ���ه�;��XI�]�����!��g����M�ﺘk�Mjb5��/^N����|�s�=���gd��:��ӆ���>��t��3=r=�8G+���Y��@���麾g�dw�Ja';���=���y=�[Aų�fx�َ8ښVYm��h��n���O�@;�
���u����1Y�3�{�O=����s+�6��?raӄc��C^8}�^rs�u��k��g��T��'�&��"~p����v�y��;;�����q�ӜO�u��n��ɿS	/S�n�t��eO�T+���G3�#�L�vt�D����A���f�$v[�;N�?8D��#S�-+�u�{8x�s's+�??�_�Ͼ��>p��E}��R��36���oGOn�0S�9\ԈV$p��53Pg=��z3��Ω���&�ô�L׈�v�s#��k�!"~=��'��|A��G�|#�kޏU����g�]9��ه��*|��5��u�޵aJi%����9��<N�*I�7�f�q#��C�,��>�gi��x�Y��zr�\>p���ĩ���,��u�@"������~���dO^&H`�9ߟo ��z�r%s'S'�~��~��:�@�{{�s�\Q�ep��`�~H�����k� {@5��#	�KI�����������O\:GɨV%���?׶��5;p���!���;���"x�A�!ܘW��~N����{e�#�<��;L����I&er��ۦ}�`��~�O���ˣV@g� >_B>��@B�C�߼�sŖ�_�x|�}�/Ƴ���*W_�\�"��_<����t��<9�����Z���7n���O��0\2��n��(�����.�Ӈ�i�P��A�����k�\�O���/��p�oN`���!����Cʹ��H���� C����B���Ʃt�(O߄'��q�
��~p���Y�>\����bL���;:6.u�U7q�{5U���V�?Of1�����n�|�N-8|�	ĘԽT<�61<XC𥝓��nT�;��u�����]���=��"�l�O�����c'b��!�q�l����r=�&Ѯ��pFώ�'��p���Ag�s�r��E0r�9��C��6n�Z�tk(\�nf��;2�u�v�S���8�Rs�p�u��ڼ�Wk���ɝ7m�9���;3r9��!�Iƌ��bFUCH���-W\tptf��l^����GWgr�nG�k�v�kcF�ݝ^&�px�y�ț���q�6h�6�}�9�����?����IQS�"[�j�� W;�^��r�c�4Nb�vI�g(hS���)�v��<W>�r�I�8X�&�,�h����z��{*{�9R@�,D&Y:����tp�x�����"����e���W��A.��J8��Z��/�zFNm���DE"���ί�Ef�/��i�� ��D��[1]o[���7k:�%�Z�[9�Z��ِzu��ո�+_4���D�����ĐH��iC��ݲ��[~��7p�waw�uB��j0��T��F֊�es�*㚚�V�C�m�� ]�0��AyA�2c(���$�?qZ�łp*tƁW^~�����*.�-Q/�)�#�8�m������#��d�P^�u@ FB�5���	3*�Qn��Z�����ލUS�l�� ����c\e�v�Jbss��\` �!�H�F�R�b����o�~����='EsՂ�8���jhG���T|��Sqݗs�R���,G<�&��Px�a7��8Q��`e����♩{te�&�����!ߔ~�ݙ�,�Ď�=��0;�n�Ϸ$��uC�ػ�;�����{V�UM����.T�hUس�9���[�L��=�_����x�`�:��*�I"�^F깮v&��32�a���g~�3���4�(0�H+�$I	��, �T�K������q�26x�Mw�(���i�g�yiSi^+��;^�}ν*Vj��;y<k޶b��3C�Hz��h"��b��/k-���;ٜq�}���{UҦ9�x�Zt�*�\�Yr���Rڪ~�޴	�V����0�Ι�r�f/�M���v���d��Q'9��4�%RQay��'J'��`�D������G~_
S�VY?U",Mv1&�$PQ�;�oW[�ڈ?5c�����έ��=g����'������7Y*4���7#7<7D�__���1b{�G��x1;?%�hJ	��b�>崲�R/�>�hh�O�	ued���`�yhBk��:4��Y8��(��"%��"��|�F����H�]ی������l�d,�1��i�tQy�k/u��G�[��R��Pxn����yHv&��b[#���o�e}�rf2}QDKq(�7z|$���^K)m���Get��w⍬o���,CJ�Q��T{|-����X<iwgvª��#eV��X;'�v�Of�����vgʺ 3��2��h���<�"=��L]��]{\D����H��Ŷ�6a-�RL�I�d�C��-�d	e�<�Y�)�v�$ܑ`3��Ɔ�fS��Vѱw+�&ҕ��Ȝ����l(X�\�^�!�����_�!Sf��˴�gpHd]�h��kI�<�/��m���i�{"}:p�sRtW(h� k�1ݎB�>9���Wg�bm��r.4�ns�f�1��`���$�M.({<��n|r��\��9޺P�;g�����_����_p��l�x.��뺌$1����X���"��ֶa�n{%mk��gB��������m3��fb5�#ZX����0��$cR�It��y#I.�Ы�v:�=����I�V�ݚs������.t'��dA
��.gN��ob�u�B%��$���}��ՠ�u�Z�a>F��8���靆���l�#I��*�H��H�ߝ,	)����oG�bߢ�CZ��W�I�5t�$�'��H&�28��O��N��7HL�0ru�o�O�9!P.q��ʣq�F�N�p��P]��
��\�P��V���#���K��Q�7� ������^�kﮃ�'(�l�P��Ip�rˡսf�w�rI�O3V�d��Y����Ƶ
�/���g�FX�ԅ�	a�S�:�UH�	���,�(D��ƿb��2��m�/�44�d�),<��q��#mYq���lFΖC�XY�.��pw+��ԋ��PYm��1��_F'д�Qm�[cه�t� �p��ڣ����T��l�\����2���9���ʬ�b�צ��=y\j���Q4�!�VC)
�_(ɫp�9!Z���p�a �u i���՜�^��Ä�r#f�^>!䏲��5�X��w`�����O2�}����݂t�icе���x�E-z앪��\�V�G�ҎJ�K��d�BBr;��Y��/+~��+�e�|`��Nĺ�+�pG�3i�^5��6�8ؐ!�@��^�o!<^'��]��㌐��q����o���=��Or��g/�G	ͩ�<2�]��A+m&N�"�i�;w�z��9���<S�.N���+N�yѯ+=)�B�`'�ig%��]>а���2�6��}�Q�)���*�諆�HA��xחW�c�@�te���VnjƼU(O�	j�^�v
殠�:�[�RӋ�4H��o/�+8Wj��ՃEF�X�O]�U��'Z�a1�[�m��,�{*C*ƫoN����}�]�#8��U�A�q�iuv�z��}
�Trơ��X�V��;�wj�(1'��@�{�٠]֗3��P���Vg[nKW��V�� � *��N�,��T�3�E�{�[Fc��{�\�1�v�XsWv^��춉�Ry[����v�9�E�X�
�ql�ꀑ�R��`���bڤRYݦ��^����f�'��6^b@���Y��5�˴�l��j���[�[��[F�=��3~�pu�7�t�A0�H�Ǹ>�E>�ݍt���܋]�kr6c#bݼӻ{�^�W٘��;�'��)��ׄ
�k�<� ��V�C����(�o�1e�F�:ɘ��煛5��;]��c��*�vM4���1�<�1=� ^�]eKj�\bos��I:������y�/kT�V��͸�9�Ժ�,�Z��8�V�����](A�l��:�ꮍt�Yo d�kj��l[��|���C��ˎ�b���9ò�;`v���]������*w�ٕrߖ�67&F��C:�'e�:�M0�cK�n����NZ��j�^r�2�u>G:9�֪L�F�]�`�����X_eٰY�4U���t�j(6�71o{ul��ʁ��vvD�S8E�e]��5I��X(OVe�
*Q>�Z|)Y��A*¯��R
Щ�s,f�¡'��wr�	�
+z3���S;�/J��W���G����hյL�#
�^���捎��e��'3�V��u�0 �3���w7�x�w���s7d�FX]Q��²����$�9#�cz.'�zݵnwQ��WS�[mr��l��gL�A��9Ξ8��ohʧ<n86țq�����;g��J��Y��uVf����b���z�u{+�Dظ\ �:� �ӼhC��a������y�U��`7`�͆�@�	�X�ƴ�%�_���#�V��ۂa�8q��U�y��Ս�x�=�d��t�gkF��[_��Ӿ㮱�t�ݶ�N��۶�V�Y{nƋO�
�=���s�9�k�ъ�X��8���h�q$z�8�7n�q�Gd6�A6���mR�2�v�%�9s���^�˭�Nq��Ȟ1K�(y�*�v9i%{^E�k����ֱ�Y��[m�$m���n@�x�;F�V��:�J6�II�RY��e��EF�\ݶ�tm.���%ܚ��Ԥ�V�m��o+��=T퀟ݦ����:9���ƒV�>m�<[�CӶcĜ�`7�C�r�G>�����M�9�ϝ�^�^e�v��]GY	�jN=��<m���܆t��Og�q��x�t�e$w��9N;[�=�.-`�{��U��X��4n�%b7V{j���m�v�Y�R{��g�ash�ec^�h����v�y��tb���c�[��a8�e�X�-��Gb��q���z�lgm�[��Y�\�jf8�;�c������Wcn�3([;��*-��y�[��y�z���}��p[����=OGH�����䝯Q�v܁��:��R�r����9�מ$�znv�cc�5���x�����<��O��Ev��p��s*���n�c�����p���(����n'�a��=����7crn�k-hI�ٴ���H�m�:6����;s��($����q��� ��������9.�mt nz�Y�"<��7&�f�u�UeR�N�O�s0��?��Z�B�s`[��]��q�k�.�W���Űv�%pW6�vN��~�[�,Qn���͹��o%��rz|���6*1���z᷌��V�>���7Y�vع$v�u�&u��8v[�Ň/���q��<v���9@�ms�X�����61�N[-a+u�y���0p�<�5ǦX�ں:Ő�;���)s�><��N9t�v{�[���Z�q�m�v�Fw>�q���q��s��-邓��\�O<�ayy3^�.�#�C�����]�=*�?F�l�(�5�1�
��;HOo�0�g�9�7��Q�W�g?
Tp�L��H
7�QEa��i!��T5��o��%3�ߢG���L��H�W�r�`���ٵEx�C�v`KDd1�X��Ύ�tu���=�u���ʂm���j��a:�;d�3m!�TC�� ��OA�W��z�m����r�Q��e/R6=;\:�ȤO�X��(��
i�-��8�fe
"��.���~�p�X~�o�N���N����ǳg���6b\��軺T�X�P)�b\h!S��NlaU����D��CI�>�1:�r��<W��i	�ݪ�4{��,I�:ؕO��{)7�t��E���t�:{=lnҩ$�G�N�0h��G��i(g�k��l_G#m�SI�"j�Y;�u
��ݷ7�h�9��pbW���j��4XMH���4,���e�4Ѵ;��=]u��A!�{��a��������yCɚ[�ZeE�f(�fCMc�]4A˲%w�J=�Uzx�[R��K˰k�ht��By������o\�n���!�Dw5���Oz��<�Ē�dq��U����xu,��>f�ޙ��O���ߧ�j�.��Lr�))��<L�v���Vb���՝z�w�\��� ��18�gۋ�1�����-�Wr)ō1`�.�Z�0�n{@�P}�j5�{Ӷ/;�%KH���Tkġ�[���m�d���)�rg{7�����*�x��ŕx�����C�*6�cq�vxò�M���ot����M���$eOh ���RnR;�hh�F��T�e��WR>�8�;��BM��$k����#f^u�o��Ĳ��)��w�L/����K���qu�?_���c�����Є���X���ptb����2"<j钦.ނ\E���W�,�<4�&(U.Yˁd�|`�>U~�T4Jf�G�Ək���Mt���pF>bC&J2��M� @�F� �����QĤ�fjG�j�"&=o���a�:��^;�$Ђko�S�ӊ�fUU�jb�����Ȅ���P�oA�p!�l>]� �3�ʴA���_Q;��"}qȍj���ʑ~�]MX��'&�ҍ%�J�)�`��zs��~W�0xd�V�^���l*��c�ᖰl�+)�ʹ�*�Z�tZ+�$�Ÿ`�+��`��Q�lKG3�l��[	2w��_\��a��"���k�Y�ԉ��ʮ���R2��F��̪+�-�d��I�^0�C�;�O�7�R�����N���=~ŧ.7T��lSL��� e����-��B���ö��=��ڏ�b�X��[b"�s�Lp� �F|�ҭ�*��>:`���u���(y����䎸*�^����!~�y����F�P:OÂ�|�J�tʯ^����Ű�,�J�2��ʅ��f�<V�l�Aն�+h��;nkFb��T�|Bi�7�Oo�d�xV&;�T�S����э�Jy\����V��O2.I�/���>R���Սn�l�,�#����g�٧G����������Y�M-�'� ���W��N���{;|�����2��+���D_��g�vQ�L��vT2���fc�]�zn��9���3��Kϑpk��k�ԙ�=�5�9<Ĩ�H�]F�ՈvN��>*5ɀ��ĩ�>l�iKf
�V���[[u� ;�	w�m;�ud�ư���/����h�.(ĎkT�1l�h�c$�އ`U�Ec��h�<�5#sӗR����,6�����u8��=v/7k�v���A��V$̨�������s�nƒ(�R��r���B$ae�]�RYǹ��D�y�O��N}z�\/�*^Εy��̐yk���->��#�2�.�ͼ7��@���0��u��N�C�`��4�'���8�i��d0�ln�m7��r<���ނqZ���NA�E�a
VǨ9	�Wu+�Xl���N�����q�G)ڭ��7g���ۉSwo���;27Z���P���üZJfB�d7���G1Q�b�;�*r���s�lAl�7o�9j(��H���qR��qѤ�+@�wd���9���c�+�{��l���\�8�*I.I4��պ���}��MS�φ���`2B2pY��)��bJݾ���N:1�g�w1�#��wniWL^���|�	�"F9"�:���Z�vm���`�3�F���iS�oa�HQ�stq�4��->	�����m_��;Hx��lX�^�㝉�R-_�FIj8FJ�ۛS�Q�{�-�@m!B��-JST��Z�AS�U�Ƶ�0狣���{@F3AI|:.�r�y!Z��.�r���W6�|gN��%v��[N���-��˽�F�G�r�N�A�ӑ�%,�iviʼa��
��8l��.�1ѳn�\��¸u�GN�5ts=N3ֻp-q��a=t�S;sv8 ;vZ��<�m�.K=�S�Ὧ��흑�y�ݻ�ظۣ֝8�\s��՞��L�0�`�qٻR�F%�/6���.��2v��9�'\lZ�x{a�Z�k����n=\۹�0�^�ݳ]b����ɳ�vLm���l��;Eٝ��A,��(1��p���s�^ݠ����:����;�Ƈ��m���s��k;=R*��&	r��A�x�g�a��?����=��A�-���)��A_��h����9�+��zO����!�]��PY�@�5c���
�q�[p)�a�mw��q]鴫K���=��vGE��+�8	��D�F4%;5�.b�ءH�m�]e������ͻ�=��?��L �E����,SQa��ι�#�N��k�]�i#�y*]8o�6F(<z!�:�� K�zŌ�n[c�(��I@Kn�Ir��|A0c�bQ)�i���z��S�/�T4�y��5F�/�˒��L{�]*Q'}�%x-j��t�}�ȯ	�/WU�=��:+��ό7A����p� ���8��b�-�~���u�l��a�I];�Lj*�Q>&�\bbf,2�_�K�1z^/f��<��53R#|Qij��*�<�n6��:� �jG.E������Hy�(��ul�tq��36�[d�nS���l�b������c���י��8W�+}�b���zJ�sg�Wvu�C\�ʜ�O���l���_O�Ɛ�Y5#�7u�z��w=�~��45V���B��v�7�A� 2���oy��5����OL�ը�o�·n��T����ݶ���j���nA��4#v;f�FL\��z�t��T������:�f�cE�HVn2z���:u˩�ϡ�Ɏ��D�*4��J�N9�r̂��{'z_ ��.jm�(�	��<ek�Y#�zJ#V��^>%��%i��(�� �.��$�H�
.8�9)���ܧ4�u7QO	��w.X:0F�8�4̋�V*��9�!�U�A��8�
k�ݸkME��j��Hk���r���J/
P�"M�T2%���E��M�|lX�t�8{Q��U:�P��ܸR�QM�g��]�!���Zg�����f�6H���N�+=�����������Z��Bu�&��h.ю�s�:���p��W&S��g���7�������+���s�\��N��Nkx�f�ٟ[3�c��T�����Yd���λUg8��F�Kb+�;]�Ӏ�\p������y��7�q���ɬe���=��fY�V.��(.�	�V��ؤ��j.L�9T�T���*�8�T���/A"����d�2Ԉ�D�z6بvlo�1M1M����4͛��b��>���*DT���׫WZ�6�T+��۷b-��گR�w�	)s�����~�w�]�8�􎙒��5^��I:�q[H�z[��ί%[����K��hYKq/�l�/�pg��K[�B?���G]tUd		�I�0����|氆��yM���n��`��ʖm���������8�x�-,��������n�����$.���LݙC\���k����Jg��-i�˫�D�x�^�E���ԈG0�d��g`���s�g5ֹ+n�N�Dp0>�ŕΰvQ��M컫t���r�6;/�%oͿ�ӴJ�9D;��Hc�jШ��+O�wXD~<���K�2�{ʷ��ӧ2T�*�q�����tOx����%_%����%�Yna�]n>{�܀ e����>Ȫ����Q5g��qZ�܎�ckAc��f������KxQ�A�'�pE~%Y��rbT�7���\.�>��
jck.U<�B;J��N�� 0_V�� �z샵���N��ႈL�7���_�ѱR8[������W�#�7 �L�8Q���,|jg����L.��6��d讥�7��6������V]϶ˬ�D	G�w��%��Y��ќ��k;�@�U��VZ�WbR٬�륆)+�M��A�����C%�ޢ�����<	U[^��1,��+Ų����5�ݼ�~�1G��� ���U�h1R�T����}����P�Qx����U�/��j&��c=0p��O���JNiا�-�m����n���GC�ظ.��K��Hm��������K����[Y}{L+�F�N�qv�0�1��K� vu�(ŭtْ\ dO ���>B�h��G�v��F�P�d�m�d�]���Y��*هg[�zcb @�P��`��pK� v�5ӂ��0D�{	�I�.��Fm�G�\Id���HoB�3�$�9�{*N���3��D��r�eT�[鯸p͊v�c�4*�-f]���)�#Q���K�e�;Y�sU��h��<�\�e) �3?p�����r�����]�{vs�uSo�Q��eTp��%b�f���4,�(/�%;�w�F�����;�8j��QGVe����h-e�(A#i8�q+U�$�-Urfwj!���J���m�
+���9�����Jϩ��.(h`q�Ep�3�xh�a?E�{v9�l�1O�Og�Һ&7�4+�0�{��Wh٣Yx����c<7�<�)�����8sՂbv$�4	⽴/�y�n`P�i��y��jVq���*�ͣ�]�W��.�����ݵxn�t��:��JVvr[h3��{�mr�Q�=�?���O��V̝X�6N�p�����q�E�2�y�&�wl� "[����>'�wE�O[��+˞yۍ�\nw:�K:�M�1��f%N[�'�[M<Nnf�#qڻmY��Z��y�ݚ��f�'<��PC�,�*[���@Y�v��h���I�K��:�eb�6����~������H�g�Kp����Xs�� �=;e��"��K]�է�qϫVX.Aūvg��8�DrI�����T��yba���=��PFx��4gu�y�����]��Bu=F2�4�(X��0:q��Ͼ^~�N;�O��.3r�"����tE�-Y��zA>���u-�s��Y��M�Բr����4��뭜ݢ�.��V�G��̥G�0'�6����I�%XM�X� d���F����Z�P�j_;h���7	�K'�jM� 1�h��Ό���,�yEx�����Dd�f�:�#�ke\X�v�EbFJ����"Z��	-�1.�xGyx�rq���h8)����ː��{[@��2��[�b���b�&�S{k@;ݨo��V������;�z�*�"�DY7Ų��K(�jx����Mv�q�
�nK�Y�� �B(T����|�őM�Bp�(/m���~�۵"f�=J���\#$	<!������x��Y�L�u�g���`h&��qϰo��ʩ�B�l�Sų�K�̲�k;��Gs�-V��u�t�+%�:���e;Ѥ�9=���8����_ef���8�N�^�d�`�F�YA����t�S���X"� �E:l]�d.,-c��Iuv�T��>�G�1`tXS$AF8T��q0�٠{���k�}OL5}��/0�^!�ML[B��>=���tߞV�$8����¦�p^���}��ҞX�99eH�6S��`�.��!FS�7B�����n�Z*,�e#�qGG1(&4H�}�n�D��2�w*5���gGP,���$�G��&�a@�qU��PycHߩ�|�v��:����=Ң�u�j�^� ��Й͹`TR�A��O��Z��M���C�(6�
��.)�<���������6�S�]8Gg�c��9��&�MtI�4�7"��>�}��o�&�}�I���9]�hw%�j8���	�V�|�U�{:��7ױu,ȼh�ԩ'݉8#P�d��\wy�A@�؋yL�<;z��E�Q�<M���xՂ<BŹΉ|�c��!:;Y��*H��Z�v�pC��e�S+��"�ˆ�a!Cm|G�$ԇ��yB�t���#c�^S��TPJ��)���*��.0U�Y�ĺ�m_Jɪ��u�̽�}��1��{�^7��^[�e����D����۹�P!ћ�3�4m徇H-۩u���L��J��^f��nb{�K��_Ǳ��@���.F��:]`-I���o
^QԌ]��QS4��k�We*�NӐ[�ңp���Z���{�9ق�s�$�T��ܧJ����]�E���X�a[nԦN���VP�ф�:�åMs>�D� ���b��GxɎ�jVva��ʣ��Lu���ھ�8{��(�J�V�k���rs,F��HxG��t�C�5f[�lf��s��X�Wb�D�SU�zOhqnǚܗ���,Y؀į��Y�|Z��-�yVvN�,�vu�s��wY�+�]f���-���B�yՖ�ۈ�M��,��,V`ʗ���#�uevig_K�*��ڋ��u,���ݶ7��t��It�d��C]�����Ur�ڽ����f7���@.���p��ޮ,��v��e��q��kr�*�\�7b�{PYw*�pP��vn�+�qJ�,�˜����+L�7V���4�n{#d1V6���~�~&L��3C�z�2��3r��x����u9�������:�WIڽ�[:�]�3�oV�0m�W�����y�N��ߧ>��%�SӝR�uZ:�E�)���GTױ�ڇ�4��.�!2� �rp�Øx�l�!,��άw2�+ye����}�s���?ʨU}�}��}�'�`������~�����F��p�-�Ҋ._�P��
��/��ӫ��Vhy9%� ؤ~��C��ҷ�K�Z7�UC������t"�Oή��^�2�* �9{#\�4��Dl�N9��YI�O����{[��1C$�1��ŭ�iͭ�b�qa:0(s��7U<�;A��4Xr~����åaK�h��	�`�#�Á��<t�붷V�u�>�&��.Z�K��<��##�{�%Gp�sܹ�����6C�,Z�qyE�����4MH�Y��O�p��2�[��R�{h�D\0��X��0�l�f��Y�Q�}�U�5g���i�&��H���P���K��U�oe{!hfG�\l��0���S��I<=��e��:Q���	D_�a]�ΐ�WW޿1T�4m��)���u�K�cy�:7��d���G�~�~=��dF4+��*�JI	R	0*)��C�:��r5oW}Da|u����S���K/�$I��6�FX��U^�)l�bFƂ:q�[휽��k�qt-�����c07�8���
�\�L;;�\�j����W����)��P��r�����\�����To�S�J���:���N�P@�H��e!��XO_�Eq�`��_l5gYJ{�X���0/og���R�ܢ	"��y�\t����f��>�γ�g��bɓ�D8�J&�Ok�Өeu�)6��ۛ'CۧtD,�Xru��δl"c�t+� �� �<y]��T�=���W���	�QG�\a��Y��2^� r;�A�P��mOrm-�=g�7�(Y�aCA"`$2���AY�Hd�,��%��r�LOR{��(p�~��;75e�_@�$�+m1T��T\�7yQw���+�8��٘x��|UXf�C�Z� ��(�-�.�1��uW��2 mh�q�C�"�$sJ��,#�朷\��NK[p�]d�Lq}�,����{m�Q] J&�`�$���}���M�hb�1���W�OP�C���#����@��	|�Y��!���=��L�����E8#W0� �����EA�H�b��/�A�4�[�lX'�!J���ג�O%!�^:�e�G��Q`lrG�v��T���g��-��	����eLP�����b��]��	7.��f$-|�.@ص������a���U�2�p%%�.���ϣB� ���%��8!!�앙�r�2��DF�|��>fHq���mV ���Þ��h�N����"(�ݺ���=i�u���n��Jz�n���r���%O]Vh���3l�5e��M������V�miJ�xwj^:��qp����9%sYt����V}�_�}v�_g�}<
9�{d�]]^�� ��`N����G9�t�&�Ej;��#��� V�r�L����h���SNz���sob�غv#/��jpg16�݀�3��[i�����H�\Z��bĈ�Բ�p����Hn�ɩ�o+��N��;��0:��ۤ1wa��u��0�M�__�I,�¸1��2`e���]g-���m�^��y8����=�=��,�� ���f��G�u��#j�����df����F��u{˗3ŢI�v���2CqF�i�䨪?Y�(�!�t�6­A�����f���i8jj�z��w����v�h� ������P�#eB�T	DDH��&�{(H��aw ��`O<U�6��r`Xa�XnH6%��J����sb�b�&��z;�Y&��e�����Q��p?'���0ZR��S΅��U}��M�y=Y���s�A9n��$LC$.&�"^RkD֖��W�@s�3E�#	*q��˴rKGV��B|�`�Ev�iy�s��ۮ�vg��i���j7MrA6����@$R��>��4%iIݜ�,�����w-�w�160�޺��J�T.�lE�(t��Siť�(`z�k���,��cI8�Ϊ4xц��g�|ylaC�G޷0��ҏ����;�ki�n�1���r#��M�;*MT�+-��t�GzЂ�YW�=K������HѻZ�[eY��)��1���$Q�+����j9�bԄ�5$��@��e��Ж̍89R������]�CL����3	�ScQ������F6������!�vf�z��
*���t-�%`�"�Hn�Q�#걲�b,�z'��༼� �2�>)V�HΣb��;e�\
���Y��)�{;�6����V�O�V$v�

.@ly����Vv�y�;�V�a���7����Q|��ݬ�C�/��4\��<9hx�->�n�|!�>���X��Z��V��Lf5��[���蔗�;p�؞ܺ
��i��P��&ԓl��iZ;�;����ZoI��ET�������9�+���89n�	-�nUȹ�7��P����ŌY<��Q:�X�Z,��r	@���5�]Xk�㞺0�]�F���ڠu!w�QC �Jj��a6�V/6k�a	�����U��q����Ax�IA��R7��PՌ$v|����AU:#
s:�d��m����4��N�5Ej�˫���N].Zr0�Y�v������5�]������9$�^K�OF�fm����C�q�>�ؼ�����kg;��&p���4b1gwy��o�Rlo�觅uTQҠ1���Ԉix%�;��+n��`_Y��"�ms�%Yညk�o�@�8��[%Gr�;��L>���>Hc��g�Ƃ1�$Uc����T+�����K�������H�]�Y�:�G>ͯ�0Eab�s	��%�⻡���c葵�O�/�t���*�(o��e�*i�v��uq��u��s����iv��s�1�g98��B�)��"G#�x=xhzyM,�;΢��3�,XE�v��Px�4�EYVC��[�ҝ�}��1�V�`b�\�|���p�Т�e�28�1IN�0(t���to�y1hRY��1�m��kY f��1i#n�0�3�T��7da��f��$TtMe���ȔY0W��3�B���Ʊj  ����g�f/�����J����p�m�"���~�UA�I�D���ϯ����*��Y֭��`��"#"�^�vz�F���&%�l�g#���nez+V��5WS�T ��ܜYhJ��=~d>ڿ�"ɃD9J�$g��6��:�<u�t/k0�0�ލ��������ܺ�#�5=H!_"t`n�6_:C=�tɿKy�L>�>��t�� �B�1��Y�J}���Ms٫d��D��}AM��1$v+��H��D�qe��{�[z�!rƇ���as�96�z��#�u��7o����G�]͚Ė�[s���"Y!ڔꐲsO�=c�b�,7[\x��Hv �[�rxO�H�#�\�B �e<5yk�K˪�s8D^��fyTwS��OL>;�mo
�*R ��dA������3�m�&n�[��%�{��eԹ��nl�p�FL��DS�J�Ҍ�K�%c��m��*V��{��(��p�|QK~@Č�+�x�VoU2�d�9�`�~� ����u]�f�G�2E�-��lJ��qRh������;5�Z���h,��(�J&�eț��-�9��ND�s �5x)��إ�jV�����9Y&߻X��+eqY5s*ԯxu�}�2���������X�8:�+Qxb/�F1V|c<"2��y�������~ŲM�N]��O6�p��� 1
䮛<P�]����58f���a�!P$���\���o�R�(Z�*
ء�{����╰pu"չ�G�7�޷��yJ��r�,u�"�1����w�+��}�]����h�����Q��ќK5���鱪�g]�����ٹ���\��W��v���T��U��q���r�ѫ�ޙ���M���n7W����hx�1ܻr-m�׶�<� ����^��m<Uy�Q�`��^$׺��qv�)	(�8O-[�y�y:�c�=�8��6۹��p �s�}������t]�ь6\&��;,͚�Yb[V�яmx;�c-�#؀pv�����=�;��<����]j]�E����Y,��ۣ����|un??!�W�9l	�l��Y���t�� ����)�ٲ���g�RSG�ъtx]-�M���.��w2��)�BEJ�lE���f�:I�ٱdַL$����K�g{ �GYpA�xi�-��r�`.�3�	�S*(�#Id��\�Y������qG�z�"1zw�U�5�H����?�U��A�o�\��y�AoT�ԃԍ_���4��#�R
0�q؁�k���T�-�d�ӻ�֓8^�ZT�`�o�V�ziX�-'Zd9o�S<�L0B��w�Z���3���7�<�{�B�	LKIF�Hk|y��(��Ix�,����]�l������^/��Z�5P�Ӵ�B\d�aUe�e�鹑O�-c�Lf��ÔHu��v��u6�B�)�Y�u;�
of簤b���4k��v�a�s�&M���`'X��Ġ�°E<q\("�&)��S�Uֲ�jE��,#��+���U�F�&��܉LgЦ�8�q��vW���>�v7k-_��h�F��&���J���TF��`��`�fe[��y�a���Y�s�[��c	rz��ō�~'E�Q/ �W�*�4%͚�ݽ�1��X`W�L�OJ�G:m[ϵ6L�g�uH�]`�W)x��<��s�[LtF�GCk��\�n8k�yO���^!r7��V?�9������:�B:��������T���fk�ƕ6�ًU�%ۑ'fM��hA�����ӑī�2��,?j�{+�WjyT#A{y����|��~xQ��D7��p�

�337ż�e���ʝ0��b�.�@i`R,�bW�M��$�CA'_%��"h4�6��\�|�c�Bn�L��b/1�m� 8��KF)pz���ћk�N�ٚs���FNәny��09�������Ny�6����N�r�i&n܁�x���6 �x4��pg��m�v�&(}h5�lַ�u�E�#��i.L<F�櫢=3��w��z|��V��E�_
)u�(;|1��� �fd���$�#��=RKZ�Y��9,�`-�&�jz�Xab쪀�����⇻��{t���FʽLn�����]`B$��0�A)��9
0Ia�n��8�ey|�:� ���7���=��"�X�Ӕ��ڱ�9WVL[��j�MU���;�Vn9B��q�2��[�[ؐ���7�����j��;ɺ�}f���K���}<g���(�'�p�%�
n)�vF����/��6�=�B{���dj��sD0MU��,weJIxc����D#�,����S��u��찵�F��=ɳm�H��l�{)��rՆ���1]�4G>��g"�q��=�x�Ug����t{�i�Wn��͈�t��L�R�pH��u�jn�U����Yh�_JH��#c��u�ۗk۷/�s�����"���ٿ�����a��fF�e� �?~K�eU<����a@��+��O:$L��?F	�ϵJl{��u�M-�]B�|�G�_6m�F8�H�c�8���21HāT*ڶ*�E�ÿ�E�bժ&�x(�y��J�Q&���'�#��S�]E� :�3$��F��9d&Spf��@��lGW�_3U��CPW�خ�@�P��b�{�G�������] 7|�J�h��ݼtR�4�'�Kn<I�<��}�T�ڐ^�w�Eso,+�4^-���.�M�$c�_+��}�+���Fn�xtb�	�%U=�
���{��=�P.�L=� &r_g`̴d��vț��e��g�4�HV�Ꙃ����p~AU�������#�����Ǆ��є���������>�t���|=��;�WqN\c��95,�� ���v�-�3)p����#Ww���Fa5��'mV�xٸ�����O�9��zL5�[ �b�i"�,����"�)h<�	�z*|k<���PÇGEފ����C����{�Kp�Z��S���<(�������Đ4�p�U��, Ӆ�Ȝ;��8��Ox����A��<C�{�g��+���y���~t_��ՙל�/;���\џx�ZnF�0���ӳ�ˇR	pT��R��-��ӂ��`�&�l���J�b�պ�͚~}H�*�NJ�9 �x�_V@B�"���368^���rN���ڧ[0C���Lq5��v5 q<Q�Nzu*�X7x��`݊|�扦����ZL���.-Y��� Y���!H��D�2 ��m�|�IL�C�5�e�}ϳNS�`��r�����
��x/j��<%Gpb�R6?�_{﫫�u���Wu��!~���2���E/bX�я�z�Z�Q�D��Y�Y:�W9Z&³]D�4�(��o�ѣfT�v�n����&�vU�i�R��eX��{U����O���.UQ�In�w�����/DΧv�$�Qely�nf��:#kt
�J�u��W��vbSv
.�V��
˥Y��7�Z��y�t|��[��v��t�:�����+#GNe�����W�����c��<�v��w���5#�v���=YJ��fn�4U΂�H{E ��8��%j�ɀܬ΀�<]�������5�no"0sι�Yy}����wf�WVG1OC�לƚ���]b���g	#�mL�V�q���+/q,�C��K�O��;agr솆Gf��XB0V��uxz�h[ۇ���a�[ia�����vR��G�.�����,3r�ok^o17��)�1�OL�JXf�n)|#�9�hMKe[�Q�Lw6��\^��SQ��<�\<��-�:WA�Y�U#>u�0ｦ�g��Z�)��
h����]J�;0��3��¨�n<��L��仲�/�h!� 4�7J�����g��}Ŗj�k3�mΊ����\A�vڈس�1vƤv��erέ�OQu�{˯b�Es�w�Ju�^R��eOU=˷�۹���a�rֶq[j��-p[+r����Y���c��J�#��W��T�#�/hm�/�.�Z=2�ߢ򞉛�^e���	@Pݳd4eib�+.TGwY��&1�sC�00(��Zh�i�=�: .#�'Q@�����x�р�����.��kf���̜�����v�\�kh9&�u��y�홽���U�n��F��{�����7]�SF�	H���n�d2�\ջuΌ�l;�qgtnJ�wgn��I�ۀtv�p�]1ɮ�p�n&��'f�C������bω|�7I�ֹ����ڂ-j�Ma���g�)�87��q�'��� �<��6���q�!�Y�j����η �\��.��֋keT��n��i�t�޵�=�P�K�+��[�7��3Ν�M�>Gm���q�Y��8=�Wk��e�3m@d��{q��/CO%�z�.6.#�gOm�����ڶ����eZp��cc���;���#�K�AN�됻n;s���9닷<KϮ@g�g���(�ck���pbN�s��6�4f{r�pd�6��X���w�u�8i�,�c�<N�ݬ�n���� ;/�896+��`�3�`�%�ƭ�kv���X�95;��x.|G�ݱɲ���N��O"r�R���l��D���6%$�M�������r9Tt�F�����,6���i(��#�n;g�ܺ�O>�m՝=u�\��÷S�A����>κ}����nŹ�T'T�Gds�&�+!p���x�\.��A!㓵v�q���S�N��&ඵ�Fu�u����x���[��E�!��Ü=v��c��C���Zz9ݱ���Sn��1M]t�t����`�]�v�-�n������pүK=��{ۦ�<��ݢ{k���k�u��K�ve���\���h�3�g�7G/����[�S��[�T�ۛ�������s���9��sÎ�	�mu=���YF�B��wE{Cx맣���I�C�I]���;<n��܅^�@U����yգX��nك��k\��n7\AUvݵېs��-5u�0��%�x;e�wk+���x�Q����u�h�,B&���y�.J!�S��=�#6���2d&�������0í޺�vI�ݲ.�1�W����ނ�+�s'H�..N�[ڶ;aجn�Q˟Z��^yc��V�l��ռ�Pí=���M�au%Xz�G�ps,��a��{s�'Q́�]�D�u��==^��8� �y3.�x�,r�>#����]W�7�4W��H���N�=ݺ�ؼ]U��î����lm��]n3��7C� zu��m����n�q;�Oa.'ŷcn��'�7:ɝ������dz�%�
G"��ߕ�5EaUS?�H3Б����U��C
�e��u�b6]�ktel���1L�b.�Z��3𖀛�[��>!�	�\�i���JI�����yG��xY�����n��1?m�-lz�D�z�=�5��RE�3R.�51�`S��D������G9��$�oeQk���үqL(4�J�Pg�N�
�s�2t@ ;є�ӨMq4�s^vPݦh/4HP&'�8���I�h��l
�������ӏI4��R�:N�=h�(x�mo����M���V]��Ya"���A��pm���Mb���4�&$\���(�u���ٖI���HF�ۇ���=�3=B���Ú`�E��Y ����5�8nCuMQ�8���y*Y�#}����t �:�����vq�[���[�[�=���эЯX����'NU���u�eAcBv�[����J$�4�i�,q�ub�z��ʑ����� �{��ʩ3U|&�Y9me��O�,6z�PLx�F�,96=c=�=�knH��x����X��j*lY�4�l�/;i?��,��^�LMJ�c�l֋�m:s&��8�Ʃ�vdɝ��㣬����&�r��4L�.j2@1���X�Я!�E���J�5�l[�Ƿ���w�:�2�n�Dkt(��H&$�L Wb-�����r���(X!�%���֓B�ΣYQ��mT�]��Rs%2l�<�ٌ���ii5O��<܉BQI9�[�	o��߽�Jб���S����ܱb��"#�]��#�kXWO$a�xo4������*�mTqk~�X�4Ѕd2�H�4)�'�Ĉ=��;㔥�R��@�7}J�Vp�d���֪��r��;��WR���Y�n_��03��B�e��o��MP=��]�T�*.0A�n��99��F���^2=5��\�p��=��Ů��$�i�j��7U�����C�N�^����\��̓�b˞u�==2ѥ���3U���l���$�8��.2f�^��������(O�)I�zX�mڅ��@)J{����ʺ]�j��ڧ�tQ#u]�C����-�l�<�)9�T��#*�6�RB�|[��PƼp���R�?�|��X#ᘡ����n�}tX����6o����h��U���%��0����w�<��+	X�s�٩+�7n���7;��x��x��Yr��Ĩl�S ���k�޴� a*��f8��)$ʏJ��ABðO_Hd��{��F- GF�pR��*DL��:�ow2ؕX+J�~�'Ւ��*;�b�z/�.2q��_}�Z����v�G7s�k}�T��+�{W.�Fn�=B�����Tuv�a�x��E����H,/\����Y����W���t�H��]��mZHE���m}�a�dBM/=Wܣ<&%��]x�v�h��o���P�+  �x��]�%,'�yA{uK�pAr�v���x���ۍ�oͧ������H#�U���RC�^>��pFL)�k�,�{�(�^�0�����a4ŚВ�z����v�7j3�P�4��D��Q����\�1�Ѻ�^�N���K�h���|�Rg�/�"5(���]�Yk�jľk�u�/���MPU���ge�Nq��w9�����wZ�b^֎ֱ���1�aIHrɣ�����Y���ClL�rKg2��s�D���;��5x΁���u�A�π�N)�/B./;=�B�U��}�L�"�k����]ZP x�ҕ4��\�a�x�CO�U��_K�%^��u���~5��S���D� �>�!y�<�ɦVv��Ȅ� R���\ؔJ��WRX�i��:�ޮ�lV��hƜâ���L���CI�{����e���m�B-�d*|�Qxf��]ҏGdԼ����)w�sВ�`�9�y�q�")�׾I�F-u�]�X�������NE����4�(����s����mk�Mf�o��w��>3!hW���PQCA��͍�w: �7�W@�|�8,+���1�N�z�yb�#Z�!=����0��D�(0��OY`��>�ު\9<�r�|KH���e��W��h�M��]u�0�ꃿ@�sN�P��Z�Q�F�Q��z�8�m������T�l�N�~����ܤw���>B�(����	q�~M�q�>��yc�W�>5l�������I���	��}�H���O8H�L�\��yF�u)K�{S��VC�L�Y�x��H�4d2[m�s��������U��YKثp�C{2�̹�F�7I�5aU����R%���7��큖���==y��2�[�v�i"8�b_�</T��z�|�����Z�֎�z	T+��n��v��m�k.�&��40��z�����_��6���vL7'-պ�8&x
�҂=bx��^a�����^E�N�9J{�ܮ;t���<��������=q�ۆBH�8�P͚�7ixM�ˀ�[[���9z����{%f}v�`��k��q3���+�g�	�cv��ێƓ��f8' ����F��v�] ǀE�m�;Xi�.�pwZܓ�zKsH֑��ʭԶ륂Mn��*�n��1ԎK�ڝ�w1U�tn�r�UXK2�M�e�ͺ�����hX�vWQ���d�_W�B�'���(S/���5Nw���Oݜ,=�0����o�����Z8��#
H`�L��b��B�33Y�J����lx����&�u������|��9�� 	'I�0_ad��o^*�Sڽf4�Jv�x[8DH��qì��Vr�Wx'�&����V���簩Z����U���Wy�qU�zj�'i����%4�l&�x��}n��g��Wx��`���jϳ%��Fy��\$2`X.��ꖕ�C��8֮BE}�HS�SI�n�n��K���0�@�"�|E8�cCy/r�;6����S�n��{C[x4����U�����$��Lt.��Aտ0�>KAG�)�����a�M�m&���	�Ee5���`�S8�u�F�n��۝���� *C��-Jʜm7et���.;,��"����3�=��'4o�JDL
ώz��[Md�+��Z��x�MI�R���A��[M/ܰ�o������B*YʐV�8�6��|K��7�%��������J�J�j�nf���ݜ��r���]�ҸU�<�����s]�o��D�}��?o5Zx�u�b��l�1�������7�3�E���<��~\ق8�b8r8���j|�Kvo����󌆥m�u��OcG0}�)���5�A��@�S���Y~<[H�[�h�,����=h� џ4�M"I��Tk�=�e��FJ�9S�m��kc�7�T��P���_i��lm�j�
�� Ju�]��>�X��,�#7�/��D+\A�26�U����5e+����&�N����m�dj�ϵ�����{S�AWD�x50�؍祚���6�֭��x����_��|��@�a'y�u!�
:7e0�s{v�;p�+n:�ѳq�\�
F�q�>��ŗ^���l�]y��1Q�B����:��=��HH]v����h�^S��ǿR�v�>X�$�_"O#���5#��Amh@����A���A��hl�`��O;�o�X�S$`���\���f1f�s6�]�s���Zܛ�����;�ʹn�6�IƬiLbꥢ9;�_<q̜�X2$��\��n���z�9�[�=�b��-@V�%4�l
�8Iř
d����N�dwFAwWK�juv�l��;a�G�v�r�p��4��U�4+�K/'vG�,�A,�gP���
0�=�&$�2��~)�h3~�N�
�J@�RJ-��չ�����1	��ha~o
G�w�������s\�o��Q��8��2�>��7��������^����Id��W⪭8�=�S|/�$��.�h�KO�()�Jz��h�y���f8x�8o� !QV�UTk���w��t�`��D*	��4i�q���LvY�iۙ�h����A�S�	21(p�j6!�a�if�}�#͊��F��}�˶�V�|5w�4O	o�hf�ELI��m�1W�urn�v_$�LZ��a�$%�BNA�� =K�:9ޙv2���1	0��+(Y9ѣ䰮��w���<P�L2Փ�Iݒ���l�-�	�0PH�dp`��|����^�{�*8(�a����֌��WOt������v�VzQCB�q]�M�3R������e%fρ�kA�A����>VFj]��ª͞J�+��j�D귅Z?]4Q��kO#6���&�\���K�+�4߫٦��V���kn�)����nT�����ϔʾ��+��κ=Z����� �t�kY��el�����$[�Q׷��6U��򽦻Q�p_DKay q^է����5�X�L��T���CJ�w��I�����2e����ͫ���O*���W<�!����c��J��U�4�c�N.x��kZ�;�Ѯ�ѽ�a3�h.����a�eɐ�P%�㒟aG�ǌe��ԕ�kN_���,c�EІ��g���~��*I�۰ qf��dc�`�ʪų�������1/��2�F�Q�
��V9e]C�C��O�J�F�
�30z�S5���Y��Q�\�E���!+}j#��C/���b{@v�F/y��������	��nFk���<����{�!���x�VW�f8$t��
Jo�w���y�Wo�&����~C�"x-5%��J�H�Ǖ�l��huoX���Y��i�ʴC���Ԟ�8��;���+�9Ay��<U�î`vi����<�D�Y�5�En4J1�����kށ���Zi�K;�k��Ie�e�uA A����됯��3U�w�*���ޫ�%�3�cU��U1+�!g����Uc|cv������H3�[�����^����h�j:�v�G�����,���]B$�%��܇�گ3v��w_�T�� R����V,��Lv.ܪt�g�u{h�<�ه�q�GpivjIQvƈ��Q�������Y[^y�Ѥx���^w��G/=[=��'^������EP[�S8��v��lqq�l����c<Ko9qLGY{ee�Mq�=w��k����n��l��H6�0�ss�7l[��i����sy6��=�7]an]�{+��lڻoC8%��EtƱ=��e���4v�v��<�sc���a��l��"�q�����:l�:�e�Kdr�Oڣ+�}���!����K��,yy:�6�ޡ���R���7�&�N}H���:
@���
��-�ʫ���ar\0:�per�Y6o3��,'��(#��gExa(uA�Zًz>��ܪ�����0�|F( �10܂��5ә	}������B�#���ʯ���É�~n��Gޗ;T�VkX��)�U^q�-}�3��2�p��!M���Y	|&�$�̎$���g��T�cC�kn���t�Q�8� ����U|��1U`<�|�OWqѝо�4q@�V,p{����AFH.E^>��چF��;n���ծ����k�}������`�W9�
Wfpv2dW*s6E����,*ZF��*|�V�X	�m,�gvxЮ�+�tg�nb��2�Bfŋ��ɷ,!��$�#�v�p\��;X��c�Q���0r�ȡ�g���\;����;�b��U�(��B���Vkۑ����ُB�V'�N�I��7��F�X_�>j�=wzF��炮�l���Vەy����[�Zh�m`<��ڙ���n�V�족��zq;�&�Ev�A��ֹ%�饪��e����ڊ���n��4�͹ι�H�fbl ��M�.U`�M^��gA�z�%�Ɓ�ߵ�EKh�л	ng�	�$w��2�1e.#m��� �̢��j9)]��$j>*��Q��'��w�S�6v����)�DK��I8,Yn�T�ٹ��Y=���a� �Ho��(���5�!��9L�ի|OυW��	�C�U݉����Ȣ-.L�UK��-�`!��q�8-|�v_��y#��>҇����e���a�v�:��me���I/b�"�n�g���^�CD�������?��mǉϫ��)���r�]����Zպ��=���dv��y�\g��Y�㌭�������z'��I�:����}�\���e���L��w{ɂl����CKEp*��'#�DSr)mtJ�5��B����@����k����,��x_���S����U�
C�i��l2~ڠ���5Y Y8!��8��E�`�#�����e��Ub��XbA�EEM��i�i�
����l�Xs�F�s�֑�18�W�Y�/�$
�~U�\�=S�P�Ȫj�z����8t_gw��U}4v�7w��8�w#ެU�ӂY���.�Ǯ�7�� t䥔'zM$C9i�D2v-�����q	�Ң�+�X�Mh�af�mc�f3æ�t#ݬ{�W!�[���`���gx���r��j_|�ecEѨkޫ�UW�Z��S��W�;���w��R���,�K�ٚ�4ocd�왏��!�J�5����� ��Z�WWmA��]ܡ��K ˃o*FZ�Ob��k-�ֻ"�Y�'G�,u:�Ϗa?V)����7k.-c#��=,���l���:ż���e�/+/s��ٓ��yȜ/1�ێ��à;elخ�W�����ŋ6��澼;]v��gd�����"]���D_]�8��l*UݢgF���gt�-���w#�}w���C﷧}�SɪvKP+�k����U�\uopN�������V����Daõp���`ؾ���=Y�3W]���å�s��8�w��,��Rf�{iF�G�B�����K�$�q�,\�
JJU��KA�k�\��i��v�Bn���i�sXP����J�=	rS0��[�[:��hvp�V+�c˭6!��o	7��l�����7�,��{/̕��2��˷���gپ�|]����N�oA�����dk�n��t���tC���[��\��
K���8�}CVf����pK�;�  ��B��F �FS-��7�U�h��00&�O>=�����w-�����g��V�D%hC$F�[$���*h�P����ݤ#�n�;��?l�q���X"̕�O���Ü�y����0oe�[+4���}�yBZ�G�K�<5��
����żh׾@r�s��u&�j�h^�5���<'���t�|�j�8�K��'���8BV7o�q�����_��C�J�{�	�d��(�nvy��;s�gL��@`����|v�uk���7�h�FL$�LD�,�%��do~�R��꒮�K�:8���{���i���X�㶍Z����[
8�0�kQ���v�YZU+�;� �fF�A�|��y�'����������	�Oc��.���Է5g��BE#�4�*�ޖ>b�"u�&��q᧣�EjR�9�� �¾nq�G��]��������!H.�s�͇�DOF�ڙƤq�,]��'@1ĳ:g+�<l������=�2�G��3R�Fz���W	{��ayw5*>0�G�S��ӱW�Y�������0+��,r��ڝ��6�D��XyM���/l�ͅ���J�q�!��錃�~��g�ܫ&����B'ҭ�����vA����CpZ|k8����S�Z �؈��ƛy"���m��Cr;��M&;k�VL�fT���Y5�⾌��E�Z���mӭ����	ԖON�������Ve���^6E���h�L$)~	H$�)%]s���bj9kq��[�w����7	�����_s(�Р���*&wƙ���Z����cElܑl�RGVk�zv��RN��b��{���"toH�y�`�@�U�
������J���ˉ��A3&�ev�S �Ϧp�4�	���;�f�&��L�1r��8`�I���dx�67�s�L�Y�:�$l�Av?1��,E�4J&Tpݑ�ǔp���n֣.y`�����5�j�GA>u�;���M�U����O����>���恙�����$��xG<����eq����j���o�'w'i�>;���fh����X��/���B�Z�oU'�9�jo^�6��"YEG|�,��V}�S�I|Gv:���i�T�ܷX�S��D�rE�r����`�w�k126����fx�������OT��S,��C/��v�ڎ���{�m݅[8FU^f�X7�;\QC�g;��<H�T���5�_S[6�i;��C�e�x�H&H�%��z�,��.�䱎x˭��qԂY�E֧��C�5g���#��=�;(a}����G��$�����ю�u�h�A�g���q��z��	��ɝ<Y�cr�B}�8�����t�l�5�bܩ�J;��7����/�m��[��Ɏ�2��;]n������,���N���iN�v�b�c�bg��]^��#u�]s���m������v����*�U�=���I����#wl��땻F��PXw�JO�R�^Nj���4��+<ruҥ�۸'Z�,�Gp�ޕ8���f��ö��!s� P�p�Ě�\F���<	��[����}�V��X���g��r��d��&5Z�U5u�+�9p#k�.<g�bth���r)r7���u�"5�UF������p!�ǁy�D]z�;�ǅ������d�ZpI��uM&�y'l; �g@�G�1[��4���O�r)ԥ������p`-1p��@/]�/)@����B�p	o`W��0?&�N��e��]Ӥ`e>\*�i> Yo�_t(�`e6D�E�P��ѓ.�]��+IG�����q�T�{]P"/J����2�k3�	��EqI;P�P!���4;��9Mf|�"k����<Kl����m�R�Q���cru ���N�I!-8��>6G�8���A�`i�j�Ȇt�.��F�ܞ2�v��T�R}��N�p��X�
��_��Q�[<6�Z��JQ�B!)
ఒ~|ޥEON�w�M�I��ݽ�|N���[�%�z�lĦ��7�۪:3bL&��{]J��&��d��{ݘl�ה�\���D��E�J�!��]a� #Μ�z��e�b���Sq���[��a������+�*�>��#��\-)eHk�\t¢��s�g����A�ٝ½�b�@���9�h^ֈ�ϋ$�O����V#(�v��jb���ZQ���)ϸ�#�/j���9�V
�ˤx�$a�����mx�cV�����o�K��܃�вo�x5��)���O����Ў��jd' �+�[~L���/qX{���¦e
^��{=3�j�p�61/�ӫ*�Z5���GOpD��g�Jg�'� ��
u�V&Sp ��i(b1B���î�X�3�R�.��=��%20ŧ��D"�
"	0�#CrI|��L#'_��`�iU("�}ݑ���~�,�6r�p�Ԅ���{�҅�0�����.�N��}��2Icm�Ar+��۠��U�W>��������{|������t۫�6a�L�²���s0���@����ŀ���o�ɕeT|}hQ@����SD������$K�°B(h+�4-�C���7�^�k$]�ᔜ�����u�ux��a�b�D� �����w[��(�5Bkem���i�S���sW�Ք�P�ީS~�>SS��ݍ�g�J.9J�	��`#��(��/��Q��$&"dmHs�O<�k1�hkr��R�����T�6��U�RI|�a�D_�7�OkG�r8�F��GΝC�+o6g�/-��?.De|J�����9RR�K�f\f,Zv^��S�6�����]ˏNݣ~��w�W$KL/9����rv6([�[���Dl)�l;�~���S�8�Gx���[n{u&"���)s���$?BH#�[�Z��b�E]�+��1�W�.
y�y��2Y1R���s���UܓHC�4��{�FM�Zo�������b�Y�a�PQ�R!^��]j[x��������j����^�9��ȐuW���W�[�4�Ҏ$D��U!el�C��Շ�i�9K(R�Z��n���@��LI�Є�Lȫ�?\	���|i��'����%�+�w�F���H��{�NwZ���W��~L�f��ޞ�J�5���6�mEE���x��m��zM��UpW3lfgZ��������._��bR۴2G;k���"l� ��N�垅o�b��ʛ�)b��6E!��Z2A]\��:����3U��iћ*bӶ��T�N��i�Nx��T���h��w�.��/%8�ef�5@o�r�`��-CxODH�{�[AȘ�E��J�|xz�<TC���*v��t�a��;�7��I�a�D���U�nx�<_��Tcq���Z���+�d ��u�\�*u⊉��Z%�Љܑ�	���866F�4@q���m�����*��u��U
�DDəG���EG�!^����}�]L����ڃݘ&����H�KR5� i�6�H{���0��{D1SK��ߊ��y�1Hba�T��|l��0�iA��s�n�ݘ<D�t��ZX� u|�{���1�㲋`�s�})�[�C~�b��'���흱�g��	5ȝ$�S��l�:��&��U[d�&��ޮ��M}�J�e�0=�����6n�U��1"�v��p?U�~A'�pkI��!i$Y����\T��E��3E��I���t�=sM(�zv����1�a�[bpC0`�S��ӽk.�ɾ&��{R��c*�K`(��Ăl7#�xy_��0�]u�*ߛ�m�X�����ܗ��1&�z�'��lE"�{�_ ��$��>�e�M��GQ�4C����묩����]H[��,	��[@�}�0T29�(l{N�LΧvc���%j�&h��d�coo'�N�Ԗ��PV�$%�+��P�2�`.����2vz��<�iz�phy��m<:n{wZ�q'7<P� �c�:�qgX����{R.�A�.0���.�P����v]�Ņ��L�/Qi;;�te�c�����u]zȭs��p��� ɸ�g�wa��V�֪�󡷀�OW�]�F���@�v������9�:%u���7VӸ�vN�Q��M��yˠn/&�����On�C�k����N.֎��B`�棍�2�m�]pT�f�����Wf��y��a�#��kLk�qak�)=oK�.���ب��؅Woͦ�(Z"B�*@��S��T��H�|�\[��tО��R2��u2/#�x|p�(w�����Vq��\�=� D��9Xm,�qx��8�c�����P1�����Hv�g�*(0ͨv�+�x*ޘ�ab|�32XP)�)��q��b�N'� P�&s�����;e��A�>Q�l҃�]%®�^��zj�*��(�a�Pd�T[�xO2���B�0�#fӵ\0^5����u���_����0슃o�-KB]�4X��HQ�^;Z���03S�l���Y��Q�wR'�AZ��{3�q�
�h<�vHv��W� �Q���a����]q���M�h���W�j[F;�e]�	�u�hº�t��<�&��판����s�dwe�%��Z￟��8�2^�NE��d��'9��L�5�P�F�w�T�tL�P�T�y�7�-C��R;/�������HEV"�q�!DK�<�E+~>5Hr��> p�ySg�-��TwxB�q}��i8b�K .���e��鲧�ma�Y%�Bx:��ġ�:)Tw�4����Ѕd�|x���u5L��7bW�*�C���+-Ԏ��+��r3Zw��\�/v;�Ř�Da ||���)!��P���5���I�L��D�'`�b��S�P��W<h�ξt�Yp?%��̗�S��`D)�t�Q�+�ā�	�BLr
���Ƶ�p�~Ų����e�7�d�������~�)"mo�;�Cegq{b$���YZ��t���q�p�6F��������fa�����5]�!A��ǧX�m��F=��7��F��ظr3,ꀊi�޾Xb��ȥ��}����b�@�_��kN#��ȶ�Q�"�����%��] vu>b�kvD�s�-��j�ۗ�*�A�H\���v��T[J�'��j���0'���J�ދ�(S�4� ^Z�J�<�����%tȵnW��ѽ*7�a�����\�#mEm�S��~E�zj��7�"�|Cr��u��!� \O�}bh:s0���a��f�m���9Ih;�f0Y2�]9B�A�ҴF�w�1���i1NA{��7��Tܹfcz�ӔT#J���c>���	����49�:�r��y��3u�����Jy,�R��nSڕB�{fS�9���+����R;׽ճ��z��N�*�a�m����X�2��������L�\f�h)ð�\dI'�0�"U��0pT��/m{�Dm�j���*�O��8��*#y1�'�X=��$j]6� ����y��^�Ig�ž�+���+��B5�2"������
�^'��s����s cX��L��K�j�9��pW�C<0p�/�k[�ƶ�������M�Ƀ��=A�IG�"��n|l��D���y5ƌ��>�����vl]l�ݛ?!5'�K���f��5�[s��]�+M2NT����h�5�á����z��7̟(�İ����-(R�!�p�$08���.Aw�m��|�}��KꤨZ������y��ټ���|a��9Q[�f�׻ƃ~xL�+;hX�H6��)qh@DA)"C�6d\�X��֫F"$���c��F�;Ʋ�	�if�ź���K�{�:���G׏���w�ep@s��OZ1�U��	���_��[��*ZD���3��+=�+�J��V�{��X�>@��=^��*|Ƚ��q�A����=�[נ����n���k�U]�̝��FL�D�A�M�]/�iS�{]Y �%1ٱ��K���R���cv�}A�C&2��d����b#f��NӫޛT�M�o}Mx��P�>jOk��H�:�E`��'��V�r�ma͘\c�|��ՉZ7L�u	�_�*c�����Y�Sh�(�uэn-���#^��|�/WC>&�JH��D����ޞ?-Kz��0������*{��P�6��C�����M��ð��"��q4���3+�]���'��A���0J8`�y�O�7do�)�]!�r��B�;},Iɽ�qB��!J�mؾ'�c	��ni��jç�Ǡ���1nF�/`�X~��N��z�{���o��d���u3o��}��&����'y���5:�g����a#�p�����m�N���ެR�N��&��h��3O1���	0����`�E������1��A�[>����!�V������	��i�.>�u��t�B���_q�pw��u��瓙��A��\�׼����t���&N�(gn�7&:��s����h/��3��WC{���2��o��Cht����`�ie4�$<�%cܾkn,�L
<�2�H;�X{��R�t�������7.�vp�6�_D@-�s������֐{٧���p\,��BCsI/1����y����3qDm���X���:�L���y���N緈�搨�����0���������ZD��zѹ�D�N�N�"㝼�!�p<��L�]x.ţSi��OuT���;���o��1ks좲��rЦN�&��}F�nTC�F,;ٓ,*��|Z�ٓ�6C���l����6+���<�m7�Ѿ�C��x)"�w�N
Wv�֩���ֲov0�8mK5$ޕ�=]��X�\���7B�E�*a̫`ʗ�p���|�����$Y�1����T5��w���;����P{^	���  qv_e���C:���[�V���D�چ���b����M<�6kj�V��'��jJ��AW� �O%ĩ�Y@�Q�U�֋)1K�C�kk������fߐ��;Y7�]a�r	=1o�ɾ���Wg��ܚ��<�VvNOi�ث�g-����#'�����q)t4���[]���ؘ&v���﹬j��i�����-ޣ�0,��L���W�X�����Z�*QELM���{�{�-^t&���wή7}�U�h��S����dF.�����vwF�sEZ֔���.٣��˱�y�ֈ�vփ6�ݽ&b�����i� ^�t�;Y��{��ﾋ�DR�qz�ۗ�4=�<�{Oj1�\H.�g�����z�
3�)%֐$$���<k��{k������H90Z;.�p�h�PX][��t��Kz4m�d��s����\-+���e۶�)�vx�Yu���m�9ƒk��AQ8.�ݏkv�����qI�ˆ�q�7*�;�pIs�g�˭�A��.�4��GEKGf$���ٮz��c�s���u��%�]��㍫F���
�:-��e��Dr��]�jl�������a��4�4x��nSx�Wm��8ĸ5r��X|��ۡ�G`�����v]���w�i�O!oN�v�ڵ��ώضLnb�u�<��}��ZC����7�k��ڔ�lyv�F�r���mQii6:rp��Om*��v,��w;�W�Q;�N�����nl<<Wa��l��K0]��\Nⲻ۞seW� �|Zy�a��\P6܄e�Q��v��s6���@��>�|a�9�����Ů�f�\u�0GK�����G�8�;��=u��$���.���F��{v+�8�
MV�*W%t�d�Xi�s��Z��Հݕ7;uV�<ZÞ�|���4�����=��㞄��s[gU�gn')M�F}`�y��ֵcKqYf�v"3WX$+9���[.c�=�]n�6�A�]v��p85+�q��o��×]��©�|�pܙ^�:hݥ��Ȱjیh2[ۗC�]��N^%1�n���e�Hl�X5�#��;�x<.��D��+�˷�*9AAv�;�ڸ@�s�nm���}k�v�smƑ���Mי�C�J�9�),�1��umc8�]����qø:�x��(9�g�ں��ktlk���'�!H��]�]s��ù��[��pss�6ڻ+k@�cY���ݹ�Q�A��Ns�m�=n��e�����&��6�[���P많*S�l/n8}�S���������݇�Y{ux�/k�Uv���<��1��濸�����r�Ӭ���(8���99b��z�\�V�och؅�kt��ӷ/��`P�ݣ��y�zV�;=�:�E���v�l���\��W\���n,c��u���ǣ��q���cj��v�b(��Y���:�k˱f�P�>��7��b�y4�����f�5q��nn�^��4�m�����x^cNͶ�]�SW�8Må�.grܚ������q�;`z׌Uts�P׷�����^v�y�ų*P����x��'�p{0�)()�Q�?�Z�b0M{�Zt�8{���Н�M�m��V���'�Q+��@��ab�đ��}3�^�ӯKC� �� J2����Y�c�Y�ݪD����:����Aפֿy�6���x����<{��'���\.�Vß6���؂�����~�����?\1c^Ǘ������O�u)�VZ��;�F��J��z$.�y��X�'ycgQdA �I�`{G�y�]DJ�[���u��׆׳ֻ����t��ׯ�6|�s��]v�O.6�{��n�S���q���"�0 �IȺ笇/FԿa�wHg��ـ��*�	&��}u�X<Fm����D�_l�f�<���Þ������ߟ��7^_�����e֭��Ԡg�1���4x^x�V�(x���z��p\Px�������K�A1Z%e�Cα��_������~�K�.K��v�\j�T��@�����VC61}�z��'��H���H9��Ěz�VN��H֡����)��9=8��f��a(f�9��a.��E�_W,�j��Ρ*X����i[��&�G=<�U:kL����"�_��]��N�Y�;�E�I|r����p���b^�W]ށl�Oph B���˔�WeFҲ�9�}�$����iN�<�~���Ou�H�Z7��+��5~C���&�ȣS�!m�"���zIZ��Q6�i�Z�-bw���˩�Y�`�[[F��b���x�͋�W�7����
�S66��4@ath�9g��c��i��6���z��>��K��TM�`��.֩�o��Ǳ��sƯ-O>�bc����o�����?h���˻^P[�;p�xm{��^���<�k�B���e��)(���/��iT�M��s8����A�6T��h��Ef9���G;�{>"���%��O�@�3&�x��*s>�e�[A��v4EՇB���G�*�u���R��f	�Xgy�lߨ��@Hdv�E�9����Z�/�Q�IR+:����8{��9Mu��ŀ���b�ׇ��K�K�2��'�\Uۿ��O�睒��-S"�k�F�V�H����	���=����,K��Z��ݰ�dc�?]q��y���̝{\۰I�t�(�f^��q��3x��6�
��k4ӋX⢴ֲ�r�=]�հ�V ��.Ժ��In�[#>� V� ��)0FJ�*�s��k������!�:pb���ghf|��.zmŘ-|�p���/���(�U��5���X:�Dn�9�1=�=�����N�HC��Y�C��5����(.k���~O|w~���}U���f����y^ۄҋ6vii�.��^��
�4V��=}�BA��LH��_�����X.:6�Hq�� 7mp��xF%�k�bx4�������V�]o�C�#�/COђ�J���jȣ��*os��6�P�<���.O_#��E�8�Y5V�|[/l9]�UY<*��ݏR$�����ȑ�<��˹�����si�Q����t�]p'�[��t:{'�#4����e2�ƒOP]�J�ޝ�NZ��r�+���I��;�E���s.�ݺ�0VN�����ַ�:}\�z�s�oj�D��E�fP���)�`�P�K���B�3�R����6;�������0h��.���x����s���x�e�#C�B\� v�v4�쩣����uHi��t��g]�:� �p���҅�z/c,W.��Uq���C�����qq_o�V����-yytxs_^�kT0�B�A�������CQ�$r$��z�1\�׻}�<�C��*��Hu��ƅŒ�a*N�N,;�-]L�[�����罐��ID�T���K�m�d�Ӱ׋�G� �}ڨu��Ei����fW~8~g}�O�D��T��D�a�,�4(�̭�x�.���X>�!�7�h�� v��)�C�:b����X��%�'ީ<�ͽ���6Ծ�MwS�8��ƐQbR8��wܫ�t���%�sH��	����g_U��j�m�._�y�䮸˹�t��io-�Yq{b:��3ZV�e��U�'2�Y��1bu��T5�����T�a�H���ࣚڙ�nT�u7�]_�+�6�\�Nōӵ;�ѵ��3�V�N�m�uq�R⸮����O9K�l�'�2v�����FT�e�X$Z���6nݡK�b*�ඌ�6��a�7lg��2;��}z��
��*���+�����t���-uc/�<��'�X����G���]9�i�Z3��Ssv��nx*ƞ��s����ޢ�[��c6�]Mǟ'Z1s�ζ�yn����u��|aD��k;<�F1t�lxw`Mb�ms����wػn���ڛ�4�n�~My�*����o�}�"�NA�1#0��Uɘ��b�ɂ�|2��b�^�I����s���[� FB�$��x^�4זNj5�o/��cd4�}�����)�a�W����B�<����fZ\E�Ǉ�����D́I�Y$q��R���{y=ml�ӑǜ�z#��T�b�FԱby��O�{zDE��L��p�P�t��9��O��%�{Ό�V�k��4!�o�)˻�م�B�ŧ���.%�wV�n۝+%w�_4�r% ��|7�����4��[��P�j���&��K6h1.�9ogs3N���ؚ.,�Ǎ�N:f����~%l�ц��[��û{K����G*�'6�9��lFD-�ő�#R-�=��2�ګ��;�d�)��h�jt&إ�+�t��r��7���;�}&�+��D<d�d. �p�����|�z���PU/kn��t�u�*��׌�k����X�X;a��`���L�`�g�5*4�����k�ZS����������q&�'vVGjHc�����cIw�.4�Ō]	��ͼ������Hi�E"�"Jx���g����M4C_]�}m��ծ��<��6w�<~|��h
�ܽ%�_M��<T���p�d��{U�Υ\����=g�Z��be�5��K��~�f9�Hǚ\��٤�C��Z��4=x�Yʫ$�_"�?9Q�|K��XϔX�~�Pѡ�g fԡ���'&���HJH��v��έ'��@ff�e�}v�;��}����i]����;Wϗ�І�lg'\Z��Ѻt��'m���n�pd����$G�R8��V�鉢)��^�Y�|��:�)^�pt�-��N����Jt�q����خ�M���n�
�����y�z�OP3ݳ������Nj�i''��3C8�8ok��;�]*w�˿-Y�i�J��Ծ��@��$��5�S��zb1����Y�^"��{>�h����;zb͗z����v`m��5�v�gX���xd2Dt0����x�
"����dZi)1a�ںŚ�����6�TU�[�?w�ܷ?_�g׊
�:�"m8�A�$T85ds��Mx
��>HB˴�����D�/��l���)iƎ�oU���
V��kp]GE�mP���ńLm��46/������
��v2���SCq�α�zE~[�����\_q\���d�`�d
���;���W��z=��S�+n�{lv'�w�vGV�܃y��b��C���oMir�����I�?���oFE�����BS����<�Eь�t���F/�����+i����{87}�93�JFQ!$�U���b�k�ϔ>�M��.�2��}w�YW.�5%Z�\�|�=S�[�U�R�;���"�E���F���׾L�ΆCM����a�J)�p:��6տ���mCޛ0��K�v)�@��N������,����+��������8ۚY�cYy��WK5�H��cAM��5`�}]�ջ��Fh0���%�*#yѻ�ASGWp�u{�*�R|Y۝9'��4"�}�U�\+jJjV��놽��2L�+}��c�W����DLe
��oט����P���,Da�������Z�K�4�*�u2�)�2$J��*ㄅt{U�Ot	��V�*��Dd�;<96γ�k�{-ױn��Y�m��E�����v��
c�����8�Q����S�y�I9��0��a�>kZ�*ѩ�coӵN�@�;�닂+�6L^�d�%I{�UW��Wo@a�~nL�c��5�+z�V�����Qm�lMl��Wc�Q`5VrYцYw��j�r�	.n��^�cF�8�\n9����L�Q*徾{Yz�m���u�°A��]�;}�,H�	H�"0��'�u��k}9�sx1a�g�zӉ�Փ�*�cH�3�^�	wG���=�MQ�C�=��-����q(a�:��_5��n�vm��[pQ�w����v�M�f����z�W�������}E�\6LP�A�o��.qf��x���]t�	��ܦJ����Ԙ�~d�\�UŹf�-R�z4�T��;q��U@�w�pթ/V�\ݯC������β7]��,\y��y��\뫊�sl�"����,���5������v�p��Ҧ���f3��v���r�Sv�K��6�NN�����xw��sݜ7��Cttچ�����k�{< Wc���(C�k��k�/nݱq��6H���%v����U���^y;m��+w/��6��:���fף��-���9��7U�t�%��W��۴�v����m�=�����hAQ-��nC�ܑ����įԺf k��)vu`�/p<�]�@Pt�:v�0�v�]�u���͵yu�0�$�M�����;�7�{9���S�͔�g�[��]�#Aض�9��,©�?0*���>�4 �1����]	#JA�V*�;W�U�G�Dgc��Y�%L&\:���XVD�7G4Z���=�=X+�򋳆��5q�#MŃ�MXΌf��Ҏ�-�(n5�;V���U�����"�}u�n�2f�&�Y�����o�S�D�\��46��z��.U镹�Y��6b�3�＇����Hp�0S�0��Mup�2��p-� [i�Z��;\�϶�̮��l:� ��qΉ�Vt���#�i��p��ĵ�~���o�e��2�t �I�	�Lt:��u|��8D�_yy��1(�u���g�ѱ\��c*q#|9 �u����z���Ѯ����XSHeJ6�G�gE�:��f��1���[Z@�;�֞�j�T�U�Z&nJץ���Ќ�b{8�X��t;�;�}7z�����g���=OXl]���y��>d���$-2��
�ٖ���K�Z�X,��n�^�r�I��T�3�����A5ds�7���`��hO�ʾ? V��F�?�g]����^�{5qX�uV�13��xG�k�c(>���&��l��8?1�ئ�k%c)6�N'
�.��p9h`�vj41����B71_f�/w7>"vuK����T�	t���r�F<��VAT2��=%-x2���~1�D�#� �:5���M��t<v�Įո;g�7Vv�н��P��س��
R/�����g����S����Oq�9�r�잿6:7�NE%�>��R�3{�XCЈc(�e7�����z�Ա��`�m^FE� ���^�	��8G|�:�{ad*��=�ǐ�ԱC�Fyz�x�Lq2���LE��y&�X�]8�]ɸ�?}��P.ńs���2syS;�d��Zd���ӥ]� k6�T�{�D�1��j��k6Q�c�`"�\��,Ea�������9�K���Z-ǽ"�+�ۺ��9v�A��5�8�f����r`<�v}Ֆ�����!����o�KM;�����V�]wiᯍ���r�~h�����[4H'+����M��sx��f�~t�̤w��fgb;�Ty�g�QY\M�3t���1wh��9F���Srq<���U4G���3/N�;�
�*��WP_���J}���ҳ���T�d���+Wr̭ҍ�]�Gf>B�0�r�aN�;�g9#�c��w�xf��ٯr�W#�YȻrO^5;��[��:	���ڽ�K\^�o]�qΨ��f����\}��:v(]��oo�Q���O"��S�$3��zr��뵞�Cp�6!��J��oѷ�l���d�L���r�&�N�������È���[�e����q}.��`��Q����V�+SU�.�U��@N�Ҳ�W(j^����Q��|��"���Yc+�fPp:VyV>�Y$+.u�����q�}��{��єp]��y��WX�$W��xEd�:ң�[�{��Vx��C%��ͤ�VrюP+�f�ebM�4Nu��7kjV9����ܹZ�@Zip�N�_<߮ܮ��<;�ӳo��u�d��"��qEV�ݝ�1p�4��jgma�����ń�D=R�U̱+r��CƳ�<����Yթ������b>���<k�2��n��갗	��ɷ���f� "�OĶvKH�Q�/u`����p���u�W���%@x�ž2����W�Ƽ6�]kT�ف!d9�k�O�D(��F'љf3#�R2c���a�Sx�b���n{�s�0�4E|��>��_'Y�*�����F0����v�আ�
i�R��"suϖ�=�)����Ru��.�Vv�v��֞��M8��8�;_�A��W�)����B��t��=��$���OQF���.��k���bD=ލ�:�p�"�~����`��;�S�iW�W��C�~�rf�������WOa�v$6kT�v_LF3D�fR�;*k�6d~7�z{aALv���で�mH��gv0,������X�ȩ8�Y����vz��ⅴ����,��9����8OJ"����m7KL��xzo�>�t�*o�G:N��k��M5�u1���Al؝�wsɖ;�ӎ*-��mZ�{˪�f���^��raS��ܢ���l]��v�V��9B��{:h�}ʄ*�q�+�O|�V�}�R�)KKEupB�9���'��7���N��9���r��� }Z���!FM�Ď��J]��k�����'\�vOܤ��o�-��Q$�F"���r2Wq��򐽝����ۊ�띹/S����U-���}�nq�;�;R��|��R��cx9�ν���a�bݺ4Şu�D8�H<�����P��\�A��L��.���Y�F����&bu���Zvz�o>����\U:�'m�f�͆���]V�S$!�[e��>�g �n���tʂ�����o����weM��/�S�2�g�ܳ�X{�
���|���,���	�&�+gL=�.�U���E�C���I���f�H\���ÿ��6�7u�_H�`��]L��WqW0��Hـ��pW�P�ܠ=:���V�p����⺼5�8V��NgS��w�ͺ��ľAjj�]�l��&D�\!]�}S���n���m���rs�+y3�
ue��R�kT�3�y&V��t���$����
��+�nf�z�lFv:������mьԝsU\��9L�>��8�;8�=�p^9׍{u�5�ns�ϣz���r��ף�iq�Q�q���v�#��Ńv���\c�C�Ӡ�6 붹h�:�{D�z���tW��v�tM��q����vWr+��6��O��۝�!��z��p�.�库3X,
r�ǛN�����5���N뗨{tfZ��vN�aJ7��8�<˩iNu��볈-�$�	"��=pw���.�>�}p]�S[��o�5�ᗢ��3;���#�5��u�tD�1��Hb�%Hk�V{��բ��ov��؅i~���1&]�Wr�^ӊ��c���TU�OX��(���oq{6eXԙ�"���ph��o���(��ea ɋ�t֌��G{N��sc�"Sx!�F8`���j�r'��0�풇�#-I�{'��g���x��c���{mû�ڎ�O<͗lm�1H�=ѻ؋�T#�+_	��H�r{�|�.@C���p�����<s�0����wGfX�MD�r��� y:�M���ŋ�P�e���9c�W�e�#�}'�rw�X�a^�Ĝ���N����ѯf�й��F�
�b��BN/Qو�!�#d����ϫ��J��7+OrM���]��a����� -v�9L��xW�N�����k�L�#��7���LQ*����M>��I<���Q&fb�u�(kS�����9X�t	�GM�`�[��4ovr�ճU�潶0!�j��̣��?�VGEm��xB�,��27��z9����T�0��?r?4����g�}�ę��_��f�����_e!L̬a����^ݛ��^���1L���w^-�T�b=�u�W�7q�ڟg�w�vѮQw㷛J־dG�E��W.�����<�G#�a�Yb5k	v���J�^���d����D��		����;KM�vc������=�d�U\0�w�8�)+i�t�̲��wf����lK��Dq�`��~vÞˣ{Kư�ǣg��vi�5����N����y�w\�9"nx:��Z[�o�~n���?]wo�\������W�|�w�6l\�x�JY)����4�Y^�N��I�E��Q:H�(����pWu��3��\�:RU�ُ�JݶZ���W�i��xq�"c�"�bذΣ͘�B�4p���n"� �M�e�|2��g8�8�D%{����n]Z�7�נ��;j��m�g&)c��7ymuЮ{��h��f눢��(u�}�:m�O'fVوfu������&P�y&:ӂ-^���Gq�)}��0kPʮ,}DaAJI2����c�s����.-|�sU£�/v)s��i�qT���x�����:����5;�vF%���� ��"8 q"c��T�-���'�K����w���5x�l�E����U��^g�yC�g�����΀զ���OC��َxsxf��V�|gqmջu�ח��l�V�:�4���E������{�o��z�1Tۊ��7m�Ku;�yZ���s��q��Έ���u�������k\(E�	#2E����3�/�掷�Mf	���>�1_dA#�7h�����t+"O\�N��c,�q]�5�u���׫?0��S,"Z��^�N�]K��yS�G!�Kɚ�L���H�5���٪)u`���8�<�<�j����8��IJ(	��!��*�k���{뛋��p����s��,Q�o+����Vdӟ�`bR�L�6pZ'3u��˼UҙZ���_M���Led����u:cZ6P��#�ͭ��aO�R�!��&]/)�%ه��m��BL�
%��Ӳ�`L�:Yʇj��yO,�:I��0�_q����'�P�a�L�1-s�g���Ls��pF����e���&���B�E��0�F]v9�p6Ml����/;��0�Ai�bM��nu��ȉ3+k��v>s�1WG��zi2��Z&pgu�����]���m�B�Ƃ��u���!�<e�$nې�*F)�P��0u帺�`�Ȕ�7�x�g��u����5<;�W��x:;�af�딃7�2�=�ڽ�3�a� �0&�q�b����������Uy�����%�Q�\�Z��w�D��Q��=0�p��e	wi��.���XB���T�D �Fyz$�j��߸��v��:�b�u�tY.���'V�G��<;�P�����4;��"�q�D�?����0��ōt�VRjcu.�J��J��|cyw5r�Y�o@�.��ro]�C���ͭwp\��
�̹�rc�:��4��kr���ͽ�ͼa\�v�(��㴧:�`������v7�te�<<k�Oҍ5o0(K���$�$GO���^�3�3�%�ڧ�N�u�s�3�E��];\�6[^J����g=L����m�{F�u�����S�k��]EŘye���3�>0��X��L�nunI�X�=B�y���x;z��l�݆ힹ��G�j�6`\���8��l�Wm�^n��u�'n[������r�}��ō�n��{{e���Ð!7r�Hn�ґ���m�[t`�����47!�^�^of��&�&X�(k����"L?��/^J�s�͉���~�E6���i(��;W<���=���v4`<H�t0��R�N/IOo�(�#�f���ų}-V��
�Z��;5K#���t�v��cU���}K��x��[LD�B��8~UW�w�fs�՞�j{h5;9����U����%]Ы�m��6v�Bŗ�4��s��a��*2q��pW���X֬��q��5�U��
s�?,狐��`]6�ݦ�R=N��<1���f�>��צH��	Q7#�8(.�W����ꀍ�tM@��F@�U�̎�d�°Îw��1���S��oE��<������O���~;�]ɨ�#��u+���$�Bx}u^����pݮ��vغ�K`tɊ�9�t��J���d�0��M���î��}��k{yQ}W�9�`{�yd��}a�k�S��(�IB�N���Ge�������q��M�n+^��(Y��'(��;�A�*ϩ����2inZ�v�ۖ�ȑ�)n��i�2^�w7�N�1�u��xe�:�vP���M��|E��X�j+��a�Vj7J�F���*6�I�c�u�?v9O,=;X*��&8�V8J�u��]:�N�wk�畈�C����7�$ ��LDT��NZ�:7<�b�/�N����7���]؞��PG#p�.�Cɂ#��1y�����ɮ�\�oڛ�a1"T%G!�So��k��'!O�4u�����c-�������;��a�;_mn�;��#�,U��7��?�;>�OW�V����utjz�7Z�K�⭯k�nN	������(8!P���8�������w45�X;h��SP;"�;e�g�}�w`�생�����|���V�#���qAr<����]^Q���_��2bxJ��u�����C�|�����]:�|3��K@R�ɵ���Y�-��MF�R94q�_x3}��/�z�F=�ݔg��g�P�ϟ�7鹳^��l��2\Hk�Їaf5,����V�3a��+g+̇ ���ƧN�^�%�;�+������[Kk׮��4���'�#Cǩ�4��z&d�4JG�95���e"��ݢ0�n��X��Ȫ�}�h��;n��������}Ma�����ok��mLj�W�P��_H�dBӐ�<���v��*�K�#��������Cm��1p�nOC�4��k��9}f"��[D<e\K��XC>��	Iq�B#�	x�:T�<Ã8/]=�;�u�\4=��������W�e<��M�����M��S��K�:��1i���f��gZ�{�{Gg�����(�Q���a�����n*=\��]kͼ�c�ዼuͪ�q6oQ�[��\�'�鵁�"��{1��i ߍ&ՉצCX�BCB(�q%n+��kk����A��O�TY��NN���.��wmv7#�E_1/�騻���d��.��%�8E8��\��:���s��2Юm5+��c�\(����A߷�l����!���o~��Sm��b���-f���y3{��!�9����������Q[�rV{K�)M��V���E}y�=��Xͯ�WS��6Ð��,���骰/N�6ɿm,3א�N4]))�Ud��9���B�Jꫳ���Z,v��&�HG�#`5����v�L��XG�X=S^�g{Nݷ!�t��rL4������%�ê;9aV��v�~O%N��M=��O+�}/~](�y���w�7q��lj���(��I��ס*�������~]0Wm{ڏ�O��p����N�a���X�;O���T<b��E��� l1�,���:3���ǱO��P�!�d��7�D�ruJ�ƱY�3Y��0�X��ZU���קP��Il�S��)��f��,���������ѷk5�Zj/Q�{sB��x�����w�uþ�C���6��MmI+8����j�8��F�=�������� �yMo�ќ,28�yc��6��'6�xlU1w�?��?� 5��[nR�	v%��4�O�ڽ��+���%���i����ꕵ/���ݒ�]��ó�l��0s�Q�u��P�����Ϩ�kU�Z���e`��yʻ�-�ةgK�-e�<�ǭ�L��k�B��pz)r���X9���޲��"�f�
�b~iĲ��c>&���fS�+~h{����)���n�b�N��V�T�(��<�
�☫����Ůagqd���.P6�g3��|�)Q��o���Н�A��
��[�|t���JY.�wk�-?m��VB��5�Lr�Wb�{
�p��a��ܯ�X˰�u3�WZW��XDo�)�gʝ�^��Q��Q�n1.��K(;��¸c�:ݻ�Т�,]>��Xps���"}wCX����f8^X�i��:�ܦ=�n���|r��@���V��Yr��9fa�뱜���j��i�����b����o����C�_e_�+�},Nz��ә�3@�Δw�W;˻<�řO��k&c����ʶ�Z=O�Ve^�[7��3*$�Iz��\Ͱ/5�Z�&��n��^��U�s���Tg��P-�{N!��
��t�^yx$agw����Yx�M�dІ�n\{�>���,��5����{T���Yk�K={l��KX��>�^ő�g��p	r&n\\e"Qגq�]�{���n.�F(��q�vz�0�Q0�>>	Zd��q"Bq����pf���m�p@��eJ�]�=�����]��y�ev�K5;G�����X�:���z�<g��s����t�4r�`v��E��	}�ٺ+t*��w��'=�s۶�{tc�wSǞ�g�G�8�%��l���U7��lonܛw�`$I]�q��a��,vٚ�.+v=�t�w,aκ]�A���s���v���f7\r"8;=LpuӺ�v�Y�V.�����'�ڛ�4�9��Z��ּ�ʪ�q�q�t��n;vPwn��pf�c�e6 ȃ��#�����OE�k.ݧw]l�^��p�8�f���-�.���[wlm��aޗnd��◴�ۣp��)>_�s#˷C+���/c��kfx�[u�ہW7���W&�w��s��*:X�>�j�2�}�=^Ė�\�މn�{=۶◮Ůݹ��uX2����v�vc��.m�r>9R���vWc�F��PZ�k�b��d�ۣ�C���z�%�;�_m�&뱮���1f���
=c�9�rź�C�n���6G*mM�B��#º-����^���/M�a�k�y�^��p7Ŵ�8�b�s�n�9�]�[g������ӓd�5���f������qm�>�(77�:�p[u�O�m۰��h��h$緅�r������[d��x�m�gpv�����=Z۳cd�!���=On:w��n����N��6<-�q*��F7U�$j)DQ�"���v�unHú��wS�O��O1>����d�-�v�[�Z=��x��e[�W��K��z#��Ỏx�۩n[��3�ܘ�	8v�(s�ŕuc�s�Ç�al��0��|��%5�y;rznl;ic���-�;av�ƭӰ��p#��Y��΢7J�+c��g��6��Ҽ�X�[.��\�`y�=���學�6v�x�J[��t����;7���羾>��[\Q/<��V��B�O7nW][�e��7:���d�N��k��Nч��{m[/�t�; �Wk���uյ��-n{t틃�]�ǫ�\5�.۵��$Ce����vޡ�:��:���i8�ݮ�u��7����rf팜i�FlR8��n��a�1p����&�kg�W�Ȯ�����7�c]���7�I��n��.K�ͻ	�A�B6��n���6Ԙ�F��/A�W�1\J�]��7V��zѐ+~��~~��!L�ˉ���B����bnE}=-�ӫ˛��bHn_����s��ذ����F\)�	J9�~�����=�,`�5��]@�5<)��V�����_��o��!2_�E���;�X~��`�ʬ���2} #Yk�0���D�٫(�{�~�e(iU���Փ�ծen�b�/^Te�=�ι���<�==��%�F��8�`���lh��*豎��g��#^��&_�)��\G��`�fmp]��1�{;"�=B(�'��׼�^�|��C��B(�%�S<��mz�S��{3���ݼ�e��ה�,�g�(����ּZ \�0fgqf�H/|�2�P��i�>J*�=2m:�P�z��C���w��g�����^�����\|TP���Wol��u����VF�OP���f`�@MHÇu�.W&������Ԅ���&d���EO�e���z��g])o�� x�Ӿ}Ow+&�o�}�juˈ}��z�����`h+M�^�X�6ggh�@�i�P�O;�O�e���]��`}��9';��C��>�~������;���y����\ǒX�2	@���]�T�}�N��+U���5��f0���r�ծخ�wQ6�P}�LW������C�)A I��g���[.�㢱֝�l��N����t�G{L��v6��U�;ϢZX+H���M#���r�A�	��$?���DY=/�^��j5�p�4����{X�-�FV��k�/��;v��P�Q�s�]��ޫ�2�����8K�D]Zȟo�����n�9�q�j���E���w<�{���r���,��j��ۛn�w7d�.�}�����T�����oa����h�^�q��V��3)�M��ӎ��a�2��xxƋ�}��ε��
֣��Q�r+�ф�Ҏ5u� �M�w�I��t�s��Ƿ2����S}
���Cf�}�:��3�R���:}��s[�}��v�r3C��)u1tS��/��3!$��5��\�Q�i�;���$جϽ185s�xV�"Ϫ���h����ٹ��e�3Z
]�:��¥����Ac���Iû�ޥ6����ެo{ffq��w�.<����"�@��n��+����:��qL᮷��g��Y=��5�3c�{���y� �D���&fCO���V�{����[���XNdM�WMWyE⩽�\�<��о(+��!�)KSx&��b��Ō34%j>���$}2d@�AR��<s�9S��o�ܲ�0�Q��Bdq][�)ڗ~����|l4k��9��z�������b�1umW�~g?|G��Y4�wq�]ݶ�]&l�Y���=�z��vs�뚟W�r���/�t��;���d�����[S����(���~^+O����k�k2����NHT�u��mD�L3�ϼ
>�b`�R./�b4����M�d�t�p���Q T�ϲ}��	�3���9'٪��GN  ��g��7c��[����|�>h�Z(~�deč�W�����h��U�cwAV���A�?u+��U��3�P|�~��a<o%0trϻ��X�*ͣ)�Dϴ�)xD�(ʂ )�^ű[/}D�GGxm��vU�f���=�����ʃii���U<B/UG�^O��v����������[i�t(">:fX9+[U�Gjs���cv�r�����㼏78�Q«��e�k�-�ᖱ�`a}]9G�?��;#o8�r�x���`h�� Ą�ef�' v�������puF���m��|3g��3���?T8��>�X/�P����Uo�]����;�˳~�O���*o�cX%2�BaFP�����7V���ˀ���3����YT����ă2�2�z1�������s�X��/F��6����v<O�M�\>#���}> ��Z��`ᵖ�ї��g��$nm� ��E����$X3�����Q��d�nj��
x�^�xuV�I�����41���=�EW�2��M�U���z*���WT/8�'��Jg�Ǒ�� �Pl8�FTp�Jʹ}I�*��;���V�c��PO��]��N'I�d�;�6@>ő>�a������7���"J��(߮{�G�f#�B��~VZ����Z�r��_x�gl�}�IjR�u�GY����j��x�*��C�j}��}.�:��UY���^����5��ߡi�")��pV���4���~��b��>����6���[WUk���0I�s�?N��E)����zq,~8|�N�I�:"S��rxI.��.�H�&�Ue�;*m��9�㿮	8��)�<x�j��/�b8"�;$P>�������B��RP�vHj̚Vr�R�W�~�޺5muМ�[��K��e�<���K{��Z��ڷ�G�򽽃 3�`�끮�݉s���s����L�
#wh��l��$�v�P��^�H��m����5�d�]g6�۲�M�*�N���އe��[�s���6�=�L�gn����wI����8Έ
��KF�r-������ ��z�n�զ�Օ�y!m6��r���K��&㇕�2��W;<u�i%it�4�Q�Rl4��wV�kwrMlF�˹���e����}�%���?~�cX貑����P�{�;���b��	C�g�����q��e4�(/
��T�^'�WUD�&�ǣ��(��Mܐ�B�'Z/¿~z�99�x�U/��f�v^����rt_��0���-��ԑNa-&��bO���,s�˻m僘`ێ�K�`�����I�2�ٌӱj��;�y踹�IG��n�^?X���P�;`=鮃g�o��^�҇�ۮ���`�"챚G1���32L�A%&� ������}W�D��r��p��f����^�u�xP����צػ��U
���g�q�Te؅<v�"����*D/�C&<J@i�P���L�Z,T�������H�Fp ����Ι�>�N�t{�'qZ�8�e�0�~Ʊ��:3kQ�[���VL�+�Շwsߪ��_�}>)�r)!Ѐsv�����v;8ے^�\b�=��\v�rn%�b2�Q)) ��zp���{T"=u�U�&�"'�`>]�-����$m���~b��w�T9��U��B���D?X8&5-+�/N|�Þ�V�~����L��qÞ�	��ÂǾ�W z�ކt�3BA���dХ��)MWΥˮ����M0{]�5�l+��*c�cf��Ͷq��z��a���P�^��C��;�3�+�.�V�+,��#<���cل�2�Әf{�f�4�Wչ���Ҳ3{�B��Ɨ�и�	��(�Y�8O�T�Ew��up,;���f碷H�9ًz%ߕ�"etu�����U����~���~�W�Ċ�R)�`
}F9RL��Də5|kuW�϶|C�8,��`��xU�*|�R~��W8�:����5v�A3��辧.q�=�ۃل@�>&��z����ƌp�%_���l�]����+���i��K����F��R=�B�%Q���o��z�F걸��������X[��zY����a%��g�I�W]aUu�nnَ���ƍ�F;�'y�pk-��B���5>�@bqt�ŋ?K,v�a���Ti��H�f�c�Oz&�����BK^����q^yX7�'��Cũ;����[>?����f�Uw�
� I `P7$d>�Z���j��k=�O�R�Sj�%{��^4�	��'Y�^�[�3���7��zX�-W����Ӟ1hV`��!
�QQJ�"�n�}�^���d��sY�=1�+Ay��w�a�k[����o���;��"�Qʌ�#�W	#4�^�,�V�M檡)�A�B�_��z3o*�gx�aW���TR5|����N�U�x�QxU��qwTevE=�a�4ͩ)���?~�L�AB�f8/�j^e����:Y55�F`�E�R0�{�ђ</
�)7^����yޟ�S�w�w��S2X���o�D�������M	0I�����n�b[�ߖ5�y2�|w�<|C7�K��x�h�Y�B$/{t\�Y]��h��1���hN;���]�_�M<��\h��Pĥ�nG�-���r�&ؖ�{�2wO*m�z�2�<ڒ�������1��+�R�P��p��ֈ�HF;󛸫�!��C�>�y�{ѱw�ȵx9}�yXe�(�X&'�~�?`�����
��ۃ���o/F��㽧�2��Ѭ]���*w�+s�:��u]׾�����>AX[�Ez��=��Z���p�փ�<��"!4~JA~8�\�砍)߯θ��h|�M?^��|1,�d�I�ma�Y�;���$�阮�q�U��ڿN\��+2H�q� m��d~H�~�!�7ɵ&�{�|.=3���gD��~A*�%?U���2;��ާs���m�N���:i���(�J�V,:Z{譺�t��nR;lX�����v��ھF{iR9c�Ck{E<����ӊ�ؿ�2c��m(Ջ�}?iMӂ�~3S���e�T���5��<"n���t�w�΢A�w��x��U�ӈ�����j�g���/�C}ˋ�7�]:�$�m�ի��3Ѯe�E�s�����b?�u����N�5�u��	�����]=��:�n{"B��?~ў������ꮽs��J�I1�]���jQ�;ȕ�٨�^3 y�<Z��zcW������p�ZIW�JPJ�����;&0�(��n+��ڰ+����{N2��s�h�<N���>~�w� ^��Y:�hw�"������TI{^�%*
T	R/2c��˂��ƺ�VK�QGٳ9��6�1��9璯4ף���V����Z�}�si��⢳*���~��f�����@B�$�Ge'�]���n�����Dփd���QY]���G��a#��AO�F��<��ֽ=���U�f�V��m
�%~%�%�SQI_�j����ʋ�b�d��zo�iW����ЇjkW���f�4)��k��T���JkkD�Ll���zv_��x�~�`z�f����C=B��y�����=�֗X��{�y��+x�\����5�n�"`�\��n��ޛ���}P�EONk��QÄg�n�Ζ+�&�⩍S����S�$�;<�[�k�`�������F��q8���i�)�m�2nT�W��v^��nͱ�e�{Er�w��8���y�nv]�ڑXu���c'��|l;�@�$ݞ���}�콤8غr9�W&{=s�=�<8�v�Mm�q:��z����ƣi�5ZѦ�7f�JX�F3p�{[c�ho<��.H�m�J�g��F�u�62r�#���*��8�uP��\)��߾g����CIQ��7�k�_.'�]�>��3Ƈ�wLL�z*���I��>�=>D`;]�s=�^$<�#�Th�)L�"�M{��I���>o�.�y;9�A7���Z#�}����R^1�ۮ�*�N�Y#E/{�m��W��~QzBU�/�~`�E�)Ʉ�y���pԗ�9�7�zG�du.ߡ/K�z�~� ��u����w�5��F��Qg�Z��V��h���I�D (%��D�o4��_�*[������ƨHkv/!���;Я�t�J�{C/Y����c�|+�	��������T�p�+�j�t^��-��>�� �$�*fI*�R.�>:�@vwԝ����BAd��A��dD�׬kއ�<L�B�ىL��L�A#�M���T����=�^��u�b��|N<�4�B$J��j�<�����]����0q�4��&��9�mq"�H�~�y��,q�"��莄T4>�G��V��\��8=9�_���c�.M�����Gĩ�1{��5}ЈԄ��M8�~:�3�Z��}��E�{=��V��&�O��p���*9���M*���L��*5ӥ��݋Ī�7�&�Cp���N�p#M�wv�E�󐺻�lX���Ob^��
�Q�%�Z�g�G*}Fe�Nvo��٣+�a�Q_�o�Y�����AsJɄ��C��v}�N�P,�{�뻕T�X��ꯆ���25h������I�:qw����y�=_M�G���v_�C$�&JD�	�g����.���]?��߈����q~�O	��9�n�5^�
�Dz�U�c����u"u�uy���:�L`������%`Ē�����;G��3��Y�D�M!�}��}�68�_t}���6˟n���'����U����;<3rgļ�W��~��������ѹ�c�X�.�"��{m:�ݭ����Kl��5���Y�����.���{렡LI2�3��$�V�q'I�^=���R$Ӟyx�ᬆOj�PT�ڶ�;��:}�R/��I�I���w{}c����X�P"��*1w�jƹ(���Te碮<u�^��Q���ޚ�2�x�x��t�#��Me=R!6���/�����T��{\="�;�����@��F�17	N�ɬ���W��Y޽j�0�˄jD��u8��Ya	��E���^+��b��lU���G.���g��y#e]�˹��Ļ�>�U����[��)�L���U��(C@M-ŕ���k���y�ݟa綻�nqC<�;T5��d7{��m��u(��;����I���B�n�-DO=�M�J��I��"�½��ܸ�MƮ���z�Zmj^�h���Cne�w��v�';ht�8E��d�����
mQ۽[iǙ2��b�D��*��N2�ͻ�Z���&�N�g2�,�����3tث�@�����<��W�Y���и2h�P�rAGM�V]�������g=�5l�Wf����Ż�����=�=nm�n��Ģw^�7�&�R�Nf�Yiϰ3��L��Y�Z��D.}��o�/�+�g�k��u��A�VC�{�u�S(|l{D�F�f��Oa9KK+3����k#. ;��7ԅ���˔�n���@��u�(���t�B��iλ+�V�(�G{��'�-r��哮k�9�-gd��.��͖8��vg^���k2��G����dU{&ևkJVQ=pDwPͲ˧ڤP���u�K�)rֻ�'l]��<ͱ�N�:�����'O*'z��m��oP��,���hfq0�˒h�E��y]�t�;1�m��r�ղm�=ܳ����uo���\�#���1c��D�WTض�̼��k]n��;����y}��"�������F���v,WV���>R	[dY��.*�����mZ�@�G�<��xE�%ţ���p7~*�6O�ܕ��?~g�,$-&�Ys��B��S&���܂���bX�P��'s����c��z����\m�r1���,D^8���9�e�n�ᝪ~`罴(�n��%I�12	����8UI�|��uO֣�zh�=o���}�Y��s�w�~y�k2=1����Y����
��\���-Ҟ1��>�*v����/ۂ��l��u���8�{E�v,�7-y{X�9����x���ۀ��wO��!ZQ^��ۏ���x,�λs��w8��O���[��*̞�9�EzMP5���!���DU(��Z)�|�
��|+���o��F�߿-z��EZ}^�5�ʲ7�}��n1�F��޼-�аl��(�u���4�65V�y�t_���;-�����ʈ${�T� ���O��=�a~
�8�����ܸ�~�蝳bߤ�����Ģ6��Y:�N"84�Ϯ�k_������l�bl��F$qf]#���+�����4�7F%�4��iQ���t�Br��vZ�A��*��pa��]�Ҫn/_�&+X�FR��aڠl��q��È�(	J��w��Mw�x��L�1���a�{N������a�����-�˒<%#��LMB��*F~7ţ���妧�t���c�8a`�dW,�Ѯs�&��0��+��5�F�7��>���$�b;<;	�;�k����Y,c<��6]��f�[�K�9`�v�yv�-��(��X�`��(gt]��$���-����{+�|/�y�e=<���,b]:�^�}�U/�&�2�fq 16���^��4�_�q�P}>Ao�xoJ!b�)�FJ	I+�����j_U�^��ߠ 2ǤE�gx�rb�/1�i�>[�d	F}�qi���{L�<��P��:��Z:��z�-���G�`��%B�d	�Fd�&C����eN{��Lz��	2��hx����1�e�DO��OM�wj�Z0������q:�b�5���:~�y�!?�L�S(%L[v�ې|��="�f�#�[�����W�t]$<r��9��ZÚp��m_}�T��������͚��Ǆ)��,��b��*B��-Iw���T�]⽍3�{ _z���0XX,��vcI�5=^�5�GD����6���d]�D�m������`�yɲW�S����M�T�P�����w�b����n��r^;K-j��Ū��=�.���6��B�w�e;�܈C��Ƿ}0%Q�����jvksu�dη=�Y����s蘎|�8M�>�n�}�=�V��BH]$�`�CJ%�����9.p��up���"�ݻK����	۲:x���#Bq�r
��rmv�q�9����N���u�Vöw/"ľ_�<JݷFu����c]65���'q���v��c�)w�'W�]���'�[�sfx=��a��=���gWms�;���5�;0���]{/8��9�h�]��[F8����%L��+ߩ�g��]�=���C�CQ��g�*|�Z��<�W:jo����r��	�ގ��]R7��m� {�+{(k��3$���$��xl[���<&���۸��I�k�����H�[A�P�����WT�[���Y�UO��%sY��}&�FR�⟔g��m ��ā(QN��KY�j�/�/FQ0+��� o�웓�E��z�ɸ�����z0�eZc3�+�_J��ᙞG�?x���t{7�2�S$�@��e�f:=�h�� ��������qBЬ����|�gJ�xk���^#�п9b�-�3gؽlx���~�����- ��In*��vȋ��`���D�.g�gXȞ�I�F/)vMM�\�$/j5��?[軆l(��3>~�B���M׀Z��7W���QSۏ��-��%z��6g
/C���^�.wnou٦{+$%EfF��aZ����ד�G)Lq�J�^���J�x�Z��Ϣ�dQ6z�L�o�����^5�W��L��4nz�ٕ��`�K�a��,@-�Q2eI�+���0f{��y㓛�#+�,eQ�-�Db�j��a�F�Ж�n���' �#�L��Ѝ�3c-8�nK�w�<��#�����4��+�ŧ��vL붪���|r϶��i�H,v��)��#������;�c�z�O�2�&�Lɕ�̞�&�Tv�J~�3��oL*���\��p<�Ո���=��ݬ:E���΋>3Ǉ|�Y3���լtK鑈�	�>�!0)�7!�䉰����	?<�vv6��l���&����D���p�~_/d�*���n)�LlW����w��Cc�w�t�h��E��g��J��R2���r��"'�Ի<81_E@���G�"�n(��?7U���,�J��o=��La:��.�ʔa��ە�s�VC���2o����JT#E��-B�p.���6��8���}G�cD�(1�&���%�5�.�K6(��2;�ɳ�X����<{����/�<m_9���6�/D�o�F���w�F3����5�'W��v�D8��6��W�?��%����2�*��n#����D�3�-%MX��_�z*��}R�ۓ2����1!{)�(Xҵu'�����aWh?B�02����C��:<�8����8 ��L���9z���2�u�>����1�_���R�㫭U��{���$���}��
��O��;
�,��X��,��3"|�#����T/���}����+��m�]^i�8A��0A@)�`_��{h�7^�T�]���)r7��~Â|H�hïz��݉�'2:aE����{��4�>z\{������Gp#QgS�^��H߾>�?����19~J�	�(�^����R�9��w�w����6�.��}����٫��M�'h� �����w�8�I���8\WC��M�2Fdf�q��nDPy�rSѷ2vH������nz]=�ٹ�]��\�S��d�K����ﺕ�G��c3�(/o�*� Q6͌f�ϴ�Z���<�k5���yg�J�چ�e��X��L��1'u����½�P�I�o���V��F����Q�@�b���`�;��?������y��p���>ot���/V����`���*Ab�uR��ia��O�/|��>����n���	@��?9y��dZ���X��I�	T0[��W���!ɱ�c��IqE1�F�)Q9m�6��~0�i��*C��J��&�ZNׯ|��ի�&���^���d2E�W�#��=D�z�R
V`t�̠���M�[w¸�- �����g�����W&�����pei��8]Z�"ό�!.\
��@z ����K��?~����&˂8�-�d�4���+;� ϲڼ�x�=��;� ��p�}�\[�a������o�h�zn��ɜ}9�2��ޥ%��gi�P�8/�~o΍uv�)<urI3gD!�:í�v �ZQx;m�<��7�����������v٨teo�N)	�r)������l���<d>������c>��K�1b�炃k��'�è�&H�	L�V|m`\Ҍ>[S�Su��D`�/�t갢���׎�mg���ԡ�����A�Y��z�^��v<�w�Lҫ�ŕv��$����ܛ����|?#(F`�&d�������φ�g3(ɀ�&n��=j�<���{3��{ҫvO��Js�{r���w�����
����Ð2_�7�?�?H���B)~6t�5���b|}U�Ww�����i�tT"p����Iˉ���b(�w�y�0�Ls�ß���u��*����A��"(A�"37b��P
<ԏ��o�MD�� uʱ-Q�ب��v�#ܳeG�Xz�*N�.���#*�.�{�+�茎쪑�Nx���F�ِlz*�%;�oI����v��Ž��[�w-�Y��5Eh<-L����,��]÷-�k�֔$e]�!J?�*��"�@�]���z��ms����b��X��\
c])�m���z�.{N. x�����<�8�Q�m���.�`8��g��!װd�7�,�ç8����nv"��6��C�Cm�� �x���x�`�oc��솂QG��� �\^���^\�Ѫc�5vĘ�ە%�݇K��ǹ�����Z��S���/��&y�snh��Y�6v	�ثٞ��6�v�5"s���A�b�v���O�߯���f��i�u`�����tJaW��g�ɩ�Faa���[��҃��9���i8�d��S����P�x�Ċ���H�&*��S�<r̮E�H�ң��h=c(v(Kq?r,��D�D����g�wZ��3�\�X��7�L�<������F;(��������ݞS��6�d)>��U� �{8o��.<�dz���p&T��~��vu��`��m����U���������L�0ȉ� L��3�W�9ϱ�^~�;ՍT&H��:�����I�D$I�5s�����p�G���:9[�Uk�{�HV
�v��gK� ��CګW��&��>w�Շ��6�u��b�=��x]�5�8m� �~�i�������H��{�F���'��DP� ��^YM/JW�psF�C�t=�����ב)u�B�M5K��t�n��~8�_i���h�&�%�צ����xN��^tVMz��F&���ZW��T=�ı�2x_��F��6�����9c�΢���W�ǝ��ӷ�3�T��j�T�?f�d������?ٗ�\�ܺ���e<�v�T���%�O�EB�u+'�ʽ7�$����vn.0�n=@a>Qyo�H���P�GS��,�$������'���g��b�`a2z;�=�
d�EL�I$fR��NR�����N�?2��g}Y{;K{�z�C2��^��=��GX"��ɑ>��cs��EU�Q�~((�16�j+���;5�*3�D�,�k�׷TED�dD�~��]e�A�Y�Κ�ji��Am�+%����X�1��.0�=� �&PR�JrƃԲO��J������x�<�?dy*9Mz�s^������U�cY��`��{}���4�SܔWP@>��ߩ����vݍ��w�&��f)�g�͇d���1�k�uw�~����Ggƹ�{�Q��*1�+3����I�"����5lQ�3s(�{/./6��9�G�@�}����>�^�f�j�I`p��� B��$�IRkGD�
�Ev�~����L(��8�=NB^���4�����(M�I�xoxȯ_D��O��r-�0��Fh�m�*�c��#�/�)t�JT��C&ߨ����� �	�?m���p;g={�Q0){j���ܻ�͕����`r^��s3��q)x�N�z�S8ff��s��΀��,��%�~��ʦ�.�s]5*�P�y��j��9�JX�i~�1Gu*���,�Z�u����㻣z&6u;rp��-VG���S�3?]]xݝI�{���%�nʸ�����M^�{�4/�>�P$��L�>2�!��@F��g�i��`��O��`W8�������$`%ONw����/�3��O����Q]�c����v�,�$I�
%"�����A3n��,��H�<�qG
�<+Y�=%���m���\\(��B4G~��jA����E��1���Ȥ^�Uz����ɇy]w����^�tԤ_��`�,��yVהj��*�m�����%�eI	2I(e[r65d�Cy�;����מ�!��@JG�
�jzfO��>�ܚ��wPrf.������mߌ縀�B�
�@�)McU�����}�%=�"��o_�o�3�3=<�4t���Vb�n�qaz}��W�\�#�ژ��@8�B L(D�Sԣ��Н$%m
y�5:M�A^�k=� ��&1%�rc��L��K�,H^���z±/�&X-] ��z��q��=���0��W�8�ݱ5�Q�����,�4��ױ�EU�P��a]�<���f_���S�\����V6n$���_��c�O��$���_��� *u�W�E���b�<_��F��f��i��a8��6����S��c�z�o��=��߇aaD�0b���b뿟���~u׺[ �H!N��u�CnݒÖkmOg���q�[`+p&;�������gk��(F)��,x��Y�^$q#'w�X�uGM� �����!>q�=�J�p{�j)�$��5� V���02�|Ah�	0D����$G�VO�����\�r�{*�W0NY�{��5��$�c��z��6^C�{(�s����>t����uF�G���.H��!� �E!�n��?[`܎b�<<��?�E�aߟeMx�Ng	��G��
�{��4�̌�q.gyM.�5y�|g�:����L��("������ yP�|;x���#/��~;H���#%����~�Q���j ����M�'N/Y�7��פ��3��\0]\2�=��A�A�1D�qVs�B�T�F_�k����}8=˰��;;=9�<�����\`�>
q��*:>e��{�������g�?���21UTU\U�d�a�fa�fT�p�p0��0���-^��χ�4�8�\x��.dP008�4(�8%΃�ڤ�ݒ%X�%ZbP_�-�	V2	V8�&d�p00��Bt���fft'a`�a�b�&A���  �3	��a�`fɒt�8�-NG���n�_-d��3E˧3K�Y1�0�)^&U�vr�f+?;Y�~[m�ǯ�Q��qfƜ�l6m����j������_���rrmr�՜�QϨ�9�c�jƛ��������zb�J���uu4�ws���mM?h+�ɰEJ�C�I���ӯ�z���w�qC�/�sO����v:Y<���7���mV�>�T�r�揓MS�yL�c+��������������B{){Zs~�6d[�9��x1�M��k��Ɵ�j���z�O��,�b��uw?��4����m�+�ֶ�$7$�&BB4�[�Hϭ�J�L�&�$a�C$�%a*��������ܡ�4L{� R����66>K���S��>/	����+��G-<g��z������}}��Wٳ�^�����^Q݌�#���n����CO��1h�)_���}���8+���/�.�a��]��|��'��N�ڏz��r��<�z~������&N�zc'�.�$�杇]=�}?+���y�+��=FL����yS��o\������#�^��-�ڑR�c.�T�~����c��}�{L5��]�C�G^��NF�Ҏ������T���tf�j��Z1�a��֩���s�wc��%� �Ɇ 8\:2��)�����g���x~
i�:� 9 s�7t��b����*�f�n1��6{���ɰ�J��E��k����U�x̯"T�c�_h�~s�z6;K�\�>g�n~�3��?{�<i�u��z;]����h�a�xtz�N�64���k,ř����Ɯ?oe;�D���D�J�ݞGy��p6��FO���}��X�%JV�a��cC��3��{�����j�˩wRҺ�͏��t��B�e8�#�ߴٗ��lp6cM���W��k��zx0�������w����h�2�l���ׇ%��rq}n��'"T�{K�]������3�c��q�����v;à�c��S���ql�s)�ᡧƸA�x�p�
���+�F��ǂ/?:����@�^��y����/#��8��9Z�3���{\4�c۔��?{KK��v�v����"�(H9�D�