BZh91AY&SY�6(���_�rp���w� ?���b^_�                                       |       �(   @                �(
�  � TP�! �E  I@
J� �T" @
(%T��U�*B��J %*AAIE(*��$p    T  �� �� , w��f���åM�� q�6�]. b:wC�����P���:�p �ܸ�P�k\�GPE%J)(�D�� ����\�F���:���V��� ���l��/�������a���R��;����w�R��x
Y���P��<����;�;� 5O=U@R*Ax z     ;�R�$PQ�,�zsu<7B�!�wC͕Cǎ�U�N� �o)^���=F�S���#z=�������x� ^�*�e��mK�UR(P*�P*�PP�����;�mJ��� 1·�\�ǎuB����L���W=F;�P���8 G����5^7��������
�<�@)
x  = �  �r�*E �������g���j�<���W,y��x�3=@�l��\:����p�g�;׀��^��w�9�Kު����T���JPN:y��=�ü�@w����zU)͜=&�;��jUy�]�6���	�J͞�:����t�e�y�P��TT%�       tJ�*����Jbo<�Ч��Q��5(q��y��W��s��B�\<wB�l��yp<�9�]�f�R���cuB��ޑc���w��	U%A  ���U,�\3�=
y��gs���͜xX�x�p=��l
���^��C�� 㻽�T�n<�Ы�Ӈ�:y�����yaT9�J��
^ �      ;�(T:�/R��z�9Ч�P���&���o-zV k;�Z�ͮ<��y۬x-^��OQ;�b����s�UӃ�z�ŝ�ABJ(��� �n�7\�zKw���g� '�y��8y7�����׳�v��� ��xe����mW'l�X�o=ʺ�                              ��iJ�       ���J       ��R�©U ��20CM0�1?�$4�  �     z�M��Td4����4�MLLF%H# A��6�h��h����zh��O���=oe{^�����۷>�;u�����T��;�+>��U{��.!�U=����ZR�W*���>_���.�����B�*������*�y����z5s��ˮ��U埏��>���__���܆d�ə��b=�Z}2�{�|����߻�/N�}
gg�V�-�l@�K8,����w4��$��WGh`s?M�,ghFq�^��t��&���oX��i��=w-툘7q ^\����q�zI��wy�ywa�-v��Y�x3V�k�>�n./���/o^�qЦ���s�n>�|!�Wr�c�COZ�+k7�+�B=��7C��骞ŀapn�Y��/rhl�����j
�GD�ţ�������7w�����xnmE+c�z�b�p�Os�֦3@O"�fY-�T�f]��ǝnZ&d�e���|�ܽY�w*x���o:3{)��ٺKŨ�r��ƮP�x�n�}cO �7�sY0\	=�{:�A���c{/n=7��Q�]����8���Y�����G��jd-ys�#�q	0�S|[��+rH�-7��s���P��	2s�v��Qޗ�;pλ^p-���%�����5�;aK�Y;�o��c��嗬}����Q%�[$mr#zi��1��8��f���*��iI0�Nj�fh��Kf.bY��Ө/�sC��֌�7:[�Z���Kݧ(�ƈ�.�w���B�3�h��߶Y�;.p�/<V���ݤ4�,3w4�v ��V�)id��G�z�7%�[�=�.��`=��sD�#��J�ݜ�xR���j<��t^�WP/fvk� C侵g#6�s�[uځ���(��a�v^9sV�)d�R�+ �����#�y�'��w�:o{�D�����&�-n-c�fĹΎ�V�������� �Of��N�te5h[����b�]�/��e�xv1\e�Ghk�Հ�#۳j��g�i�)�9:]K��m'\��Į�r��mX�����us�n��wC��R̘���J�iշ�rNN}�I$`�(iIV���g���3�*w��� ����\�7S�ы��`��qf�6����s�{f=*ѧ�	�d�P�,cN��	���]���4e��������1TN��0v�5�I.�Z��ĺ�:�h\�KG0L�Y�j����oT��$�X42��8i��x���Doj�����v-d-���ҵ�;�n�纁��KsuZ�w���smԻ&.:ѩ�h��i�	����7Y�i����Foa�����uق7"��P3��E>y����x��Vv54�Й2�+}ؖ��;u`�Z{fږ�;�����ȵd:г���[�"��h.�yt�q�x���WH��4����a�����*+T������ƛ.�Lѝp7S��P8���:�9��Rgf�J��ë
p�_D�ɽ܍�J�F��p�x<8T{������4��;�m:�	��ihT�aۜ4��b��e4��yXH�n"w�$�M�,�~����Co#Ϯ��l��{��;DF�O$L�����vnL� ]ܹ�f�D������}��.r�����@���oX�Y�54�<�Ê|�����':f�mEyZ�<���0]8+uuO����\Ei�-�L0���e�Xh��r&�h�G\й��7^�0.}�q[�Ǡ���˩�6���vEyCw{c ���u7��G �����\����x�u7	U�1v���D�l��w	�(�e��-3l��9ODnv32w��x#;��$!A����y{�wU���vӮ��GQ�.65��^��50��{�&H�,�/��/u3,1tø�f���O=�˫7�/��,g�@V,b�"��䢜�H��tÞKD�t�j.Wg�=5P7"�bk
��գ�z#@R-9H��NoH��o��!�^ㄮ��ٿMˋ���=��q�m{n�X�7.�gK�{�X�#�u����������fk'��Fut���f�GA�;G<����2�H�n�Ci��F�+k�L&�}  \s~��Fǎ���9>a�C��ٚz�.�Q)�R�RÚ:����In�X��\�b�@��a����e�`�M�;#��c��h��e�� 7�h���� �Q�6\x8�ե|T���V���+����="��g�(��f��K��۽w�|���նL]_j*u�"Ih���qgb8�uRH�];�l��A���I5L4=��x�ɋC�z=!{�]���c"�
��d�Z:Hp���˨����XN+�ۣ@��>��WD&>�Lp��VEL*�zoM1���e�\��t�L�P���:[Cy�nw���^;��'h#�΀t�"���j�՘~��|��-�G�K%qnuy3�ѱ��Lׯ��ӱ��ʴ6�����1K�̺mcvk��۷�{x��zsg59Bv��LY*��@�6�
x־_N�{m4I)4�C�˯v���'�բ��'b�Äob�pN�w�e�|c�zՈ(J�ݦ�\;4v㱛���],y,Qp�׭=ٺ�ٹ�"��Z�͵ t�Z���q��va��L�jk.T;*�mw��kq	����:�4It[�4���!EG�̹n��Y��#���/��h�ڕ0����A<��(
�?���`n�����ƴ�`<y�w���w�WM�=�f�۸h�6v��#{����܍��M�N�djr�%:�Z	������yw�{S��r 6��S������M�"�J�Y�;��u�9�{�u��>��PU��Ñ��YN���:�E뛸��'v�z��i s4>gET���<�բ����s�}�.��$�k'DNֵ�F�rm�C�X�4�37&��8�غؕ�Fc����4�[m{�0��d����샚�"��h�sP��w�tZ�;��hn��X�!k�l�Ż��ٷ����X^���vv�7s�}�܆����PZý�WiM+�Q�zZ������*͓)���a��G"�R���ه�Q���{9��-;�e�7������J<�1�w+�vs�Cg+77��ѩd%�f�ˇo$�@���7�W��0^�8�/���ag9�w�T��.Ե0��T����8����don5Rv	�"��:�]�wdsn�a��-�s�ೋUR���\�</e�2gr��?��v��ʂ[A�l謓�7zh�Zk��)v,�����3�{.�h��j�6��U>Z8��|K���;e�NO^��������cǐUݙ&�Pאp/�s�u.X�ҥ�=�y)�O<9�a�����v����YK�<����CIx �sY��!�s..��8��}��᛺��.�w�{��u��{�ӡW��n�]����f��ޣ�)�n7G-���k����;\8�bG"5ga{�dkh�7mͩc�̵e��\G"�	��KZ��uԘŗ��gS9-��_�SL��Ӑ<Vgn�VEO��`3�˃6��U-�)6ގ�suS�x,j�A��`���)��7��`:�]l�$�WH���i���|�,@�#���v]����i� ���#�.�v��n���n��yky��	�Y��i4���I�d�K4����{����
�$���;;5���d�8cr�\/8R#��聛��U�� �7a鷛c;�1��\�9ݹ�V��ۛ�%�}n�wL ��س7+�)J)-q���0X����aCov>Ꮧr�ww3�e
�e��v���bX�����"��؇W]�^<���,>�;�����pv¯jo��˅�ed�����	���8�8,;�-ыhb�qr�վ�杳{.�$����6-�He7{��80�:4wY����&�yCx�~���#�Ȋ�X�z�?٩���wy�AzA4�o42nB��]��֖��9f�ʹ���:T{6;�Xc�/NRc�!v�M�|�乖xZ�k���3�@�CM蹽چ��W6�7�-*�n��x���+^K��=�������}�n�I����e�W��ۭ�$#B��3GQ�y\�z��q�*Y��Sf�=�.�V�n��Qǯ"���p��%kz�,@��A�:C܀�>J�;��z"8��4i:c磯d����� O{ב�'�NK{U:cE�ݹ6L�F�N��{t�Eʤ%�Np�X�L]���V��s�n\��c�~�i����ohѵr�tvT��Mw�EZq�#w"���;�]�>o:���/JaM�R�$�܍v����S^=�����vlV������;/:�{������J�h�gc�1\�ٷS�6����:�8��m�&�u܍��d��dX��׬UT�����>4s3r�&�!�6�Xyt�1@F2�s���	��9�t���yđ���$}F�5u#�y�$t7�� r|�_��6{�>�:�\���)����wy�����;�H�8�����wl�i�&G�-�:���pނ��̕��f�J�D���3�p�v��@aL�9LG���"Q��S7��E�d(<����]��ۙA�|@o���s��§g֦�nE����� P��vM�GP揻�P�?���嶖$X%�}�р
������Y�tȎDh<����w^t��\����o2�.�F�*�ݡ�m#�E¾��M����7:�k[9ú�����,'��]囹7W9��j#�6&�^�ϻ�E����VG�$�\1c���ww�˷/4=�U4�t��{^ �5Q4i�Q���.n����:\�7�ك��a�#O�.��X�����X��eD��5�+�>F,N%7#���z�:��\����Ŷh�gqxgu�v��Tg.R��,n^�4�,#&=Y�Nw�4S��,zw;�=�7�+&���*���z.��a�U��n��nۛҏ�n��_�X	�/���V��vk%Dy��dn���F�3� u��˰p�u,L�k3�i"�\=��9z�{�v����^�hNa�,����� PA`F,ݒv���jˇ� ���92b�]�wgZ�'8�VR�I'gq ^�O�n�ל��Sf�k�3P]��W.u��}l�w�*��圁]!�&����60���l��]inC�ٹ�W=T��2f�w�-;�����;������j@�q�Yژ��;{q�מR�׹�z&�[�,�|wM�1�6�X��j'-W�Ȳ��b�ͷw�LXF��;��.�훏6]=�ˏr����$�u�]��1Od�-�+��*7��*��t�Fru�sw��qX]R��ׇ�tr�֯#�6.���#��':�(��7�m��L�oD<��	���ط��ʮ�z�.��q.�t�� ��V���Ϊ�&��	S[��c��WoǦF,7���Wk���Ô��ݴ/p��8њ_E�"s�+�-�_6,J��Q', ��qwF��.@0Q�;2k+OŌ���c��l4	�H@��p�/	<�KN��{��9�v�z��U���z�
��F����!Q�(l�������γ8r�.y�9 �l�E�f�K�qc�,X]Xv��U��K�ek+���~�rby�����AȚ�ӜY�v����X�ë��C��4dz��=�o<r+��������읝y��6�O>��ڃ*��ܪ�
j��&^��+af�$oGIK�t�U��9�U�`�_*�xX�Դ����${n4:蝡p"�,ZO��E�l7�§�f�S+᝻ϸ�ǈyq�tyxz
����G��.��onZ)�����o�.#�h�(6h	7��a��u�0�{�^��nE�Lv��_��lC9�&޺�3�gl�E���#;i|�kա7��{��N�TEM���5��Ѝ'E�q��I]&-��>���ݣ:�)�ty�#�e׶��+�Y ��3��B�)[t�Tޠ�}�p�X�ۜ�2@=p�	��1�b��vo�m�6ԝǗ�}���g-ܺBC �5跎�GK�')����q�^S�.8�r$��Fkc�G�s�+�^�KxNG:kO�C/���M� 8R���$U�x�Du���@��7��WZ�h�q��e���V7*���<�����v���8��ۺ��Gul,Р}�j�F��L��7/8�{-|6ꕝ�����M�O�1;;>OqkX�$F�f	-���A�ޏg ��WI�#���z6��Y�ӻ�=Q�]Y�T섬p��.O����5���@��^�0��8��)�a��Ǻ�p� 7�}�f��:4�t��[�l#��b̔�f�s��.�۫s�;oq�y�RF�b��N�N�l��[�{V��b=kmb��;X(|�N˹�S6@z<	w��{Q/;�ˁ�L���a������溠����VP�7�� �s�ñ�M���K��˛�Z�6��I�׺�u�c�/L��q�0A�V��hJQ�<�<ŢgP�BN��c|u��qۇxo��Y;�ɩ��}��M��Dr�k�sJa�	�0Q�E�����^
m�0N�N6u��6�w��.�nL��PZ��:I�h�ƭM湝�;K��]����Z:��hF�YϯlL^�й���=�r��S�y����6�T��r�^���H���.�g�f�WY��tc�w!fv9H���{w� 4�4�ۇ]����~���3����Ax����������'h�e�� ֚x���Q��U�k�8�ƭ���{R}��Ȼ�n7cZ�Ƶ���}x'��Œ���ucaF'�6�(���u3�� _%�r�b��͙I\Lbg,�V~�<v��ue+U��ŦUM�)����_��;WiZ��^Mz�kT�O2ķ�ע�S��y�u��ohv[2�y�7^ܰ&��)^[ǒŻ�{4,gq ��쇣�Z؆U��>ln��b���؉ldM�.��x�s[7�6=\�՗������������k�?�����w���$t��Q�<������:�3zNN�s�a�m����<n�Л�E燅P�=���z��NM��ga�s���{X��2���{�Ą�����5�s��7�����X\��Z�k���v�`�۬����ַ0�x�><2��'te�Α�<`��[��Ozu��9�{c�dTB�mp�X���Ľ�(���#R�"��a��1k�ۖ�܇�zd��燥�ek�u���>n��G�'�����6�I�;;v��PL"���n.��/u7P��4��^ݛg�^}&۟b�x�"94���ƽ�ݵǲ���^�0�c���ݬy,3㱶��h+u��v��{�i��5����tavù���.�atv �lm[=$�Ͱ�kb��C��;��n���\p��=䴉�؞.lm��N��Kh��i��^0kv��zյۯdoh㍺J���u�s�Y��l�-˺3qg�E���]���R��m<��"a=��:����tx{{�����O`e�ۮY�ʜA��c���p8ٳ��I���`���C����V�T�v�z�;��e9v����'���:L�Q���w��{un������Ztn2뭴�vG\I��6X��G6,�f���W��p�r�-ڍ�vK���5������+�w9ɀ�<��gp����n��N8z��C������WV�"k����P���x���t���-Z�<��v�[��k�Fg����7G:�td28&�6݂;ny���-��lƲ�s�{G��0���c�v��y�
����d�ǲ��ez1u׀얢z���\;�8y�nlgb�4���-����;q֮3y�+��=�����{��\���p]�q�6�ܻ��v9�N�ջqO8s3�6�(z6R�p;�㗤 /7�]t��;t����Y/
�pi�㲉sў5������\�^�h�&��d�v���M�nv�n#ɩ�Ǝ7S��н[�Q�<6utc�i�lz��c^tx�{0�8��M�r�k�x�,m�o<��c�;�<޷�r����� rC�v���r�Ϭ�;'���]u�^��b��tu-�B
����(MX=PP�VԴ�q�*�*�|�Vϗ����i��������Y�����]��>#�j�F��M�糗�i�Ļ�P-v�����u�8�qm8$\H�mێ�ռ��g�WK��rmv�8<8�lpf�%�[mtv�6W���g^�����	-��O/+�Z�s�#o*F`�D�҉�JMT�]�m4m�$��a������{l����뷑;n,��k�[����rC���	֐�㭧��u��v]��q��u��a����T�5��\o^It7n�Ga��{iG��mʜB�0���k��+��UO`ہd�%�7�F]�ބ1JDF6��� �8���6��%Bv�:#n��'#��nN���Ӯ����4��ש9�9죢�v�ɦ�����NN�nz.�yn%������r�&�nַa�sN�n�Hwl��t�&,n���'A��5<��훅�M����M�xwa띷av�'E]u��On�5����rCȏ��m<��7�r��].��F|ļ��c����M�����ӏ7sk@��CО{!�f��m^6���d�ۢ8��Cn~�=�̝��ڷ�xG�v�[N�#1E=���Ks�hsv��ִ����:9��p�ӻ.gu�y{G�Su[խSړ���z�0Ť6~��|}���.��p[����3�kŠ�k\R�K�&\����okts��c��z�&sD�c�gls������3�h���p�)�� /-��d��Ʈ׷<�{��.{rnt3��9���M���l�g��v.��b�n���&��s�\��ם�h��0��s�ݴ�(�/v��l�7l��x���8�Y^�'uL@Њ��`���1�UT�*�lE� �(Y=kunwVyT�ᣋ7����ꀎ����I��v�d@h���n��Ӵ`z���;ۓ�~�j�.	��j0�խ�d�6����9D�]M^xNG�{q��7��;�J��o�ɕ��|�;r��.7nx�/��vF�0·�N�����y��p�]���ޭt���n��sg��n�q�j��u����EGov1�����x����Ն���6�7���m�볧�ؗ{9���{Q�ӵm�g��>�6z|��i�!�kk��vݽ#ۓ0�^b���{��*0&f����6;c�Ҽ�;�B펺�\$�N콘䔏D<79�c;��s].��	n���8���Gq��luv��^���˓���c����h��ѣ&=nM�V3n7�d㺴��І
�����;��m���cna���j[)�����	�&666�ú�*���}����q�t𽱪����۝ϓ����#��k6��;i�1�J�G�,������g���q�\�ط-�+<��V{`����<K��F�������m��ɋ��Hw<:�V'��fț�]\(��\�{v�!K�3��{;..�i�#��S�j��Q��l���#7�rn8�^�Y�s�V��8�4��M��Ͳ�.��c�����v�]��:�Wˋdf1�^�E��͎}>7]�u�r�k`F�bۭ���-9h�S+�mI�n�ގnq͂A8
���0ʝ�A�,5@�iB��ζx;l��`�;g�eݭ����ɽf�r� VY� 4h���۪�ӍE�x��^F���ۓn)��<�7k0N�۪��|}����[��,m�v���t�!��K����듒#�=m��]d��)S[K2�G#�b��!�\������q�wg�9�)s�I�x����:<qkR�=�o�w��d�c�.��:Vt�j�*��{&��^���1Mj�[x�1�糞nw\�^;�K[��h�����a,�n�<�X��e�2�[���6h����ۂ�v���Ų������u�fXI�͊���b8�v�۝���/^㵰T�8���Vnx1�/6�i�v�l��w;���Q����.t뜻������D�@u���9غ�	�x�x݄�1�s[��.�x�]�݀�dۓ�k��Xmz��6�J۠�.]0�*��.��p'6x���]���\����f�.���d�=���y�^N�k%�ӳn�����㓗�[�,˼v���=���V��<]v�nֻ>�Ӹ�=d��ќ��K�d*�\s�\ǎ6��+v|{yT��E�<[��K��5���V�H����ۉ��z�|�j(�%���)�B��u�C��Ľ����K�͢l��卯7d��d�r*lI�o>�6�Pr�}����|�,9ɍ<��n6�b�۳�)Ǟ+�e6��z�b��5��9I{x�'ugS�qs�ax긻^^���ح��=e|���5�m�;{��;*<��(�$q���.^�)��l����9�v�x��{peXEn�n�5�s��e��Q�����v{֟ ��K�����su����	�%����۷;r
%�<�*�7���u�:Q4�i��6�q\Ԙ���04����'��_w�<u�����ݮ�cno�e��Ν�G���/.��+��_I���F�=Z�Lq�ܝ/c��(N6ş7/1�u����;���SA�ͷO�ڄ�n�]b,�v��Y�s�-�����s�uݐz�t�''3�u�狇�����A�\c���:0�Q�ws�5���J��+��N�=�wYPF'����fklb����v2����������غ�	��$[ɀC�I��\��U�uZ2�������y�k{p�=�wK��;T�E�5�H�.#^è+<��z�*c�㕭�vM��ˉqjӳ�{	ۍ�M�����oMΛ�Ui縷��6g���n2u8׻q�9..�:�v��[��=s%�F�YLa�pvw���ʕ�Hݓ�.�(=#�]�s��S�X1nz9wVB���2h"�X�[+dq-�v���;k�/G���Fȣ�ўN��<�V%�3�<��>��x�]���u����ӹ����n�ru3`%��kO�P�;(��^^��b�=;v{)��5��kM؎8�6�;k�xJ�n݃�vr�h;b��q�ΝǇh�G��u��	����֛��{�t\�����c<e�����Ќ����r�;�]���eK���A] ��m</�E�sn��]�d�ێ{I���c�]ڵƟE���3���v�;Fۯe�s������ڭ�k���A�ۨ��lm$pݵES����n+�9��n��Zx�ܝ5���r>�g�E���'��r����cӸ���kp�鶎�R�-m�"�����]����sֹ������4�t~|����0�E�>�D���� �q�l6Ǌ��'<x��mחF8���Ȑ��pZ�(��8��`�	�у�".�v��#`ɶ=[���`z��&����mihz�J�un�;^���m�P�v�«MIۑ�P�y�ź���nյ��ǋv�c�iV�7m��uӺ��n�m%�n��b�s~j��\r`�" V�B:�(��v���j�g�%z���bt.�����h���]Q��=¸�z6�v@um��ێk�۳�7���[���;
�;�n����헇��ۉ�Ҏ��n2okC��K��)��÷u�����7��٨D:T*;u[�MT�%	[e��4;Y�jsۭ���/q�PM���W(Z2U��Ǆ��t�5�)�]�'�H�z�{vG�`�K�O*���Q۱֭���x�=�_dsr<u�u�]n�h���@8�͉��^.v�g�7����λc���<�lkrBz㣎�x����dƽ�2AW,��6��qی=6G��9n�Ӊ'=��sm�p����D��9�v���]k���bz:��CCf�\�[.�ꣻ� �=������wk���G[ۮ#���R�������[�v�vv��$`����v-��<[\��]�n���N��yi˭�v6\��Bq�m�i�wnz.�x클';u�8�zs�{��G�a�b�Z�p��Ǘ�ļj���0�����n�r����a���A�9{oWn|�W M��v�����������m�ӭ�8������ۥJ�%My��+Fy��t�n�x�㫎nfl���Z2I[�n�����n�۶��ɑ�6��9|���R�W?o��~���PW/�~q}���<��߆�ww�q���s����^�:8�����=�9/�ZK�}{g@|�<"����nq��L��;��9�ד�5�}���G�v�SC޾/|�"�}|�;�ߞ>xz���B�����ޞ���{���&�s|���Lv�L�Ydk�>����o%GqX�B�W
i_oicI<�F^�B�/��t>eX�E7�\��y�!گ�=I2t~��$����;��C�=Z8����k%#�.C���H��ٻܨ=�\w}��|W>���[@�+��r�i���߫5Gu����0C�,sȼ�yh�X����̻��x�k�B�+�D9��s������_qj���N�J��i���)+��0n���`�
�ѧ�t�g����<�rR��k�?I=w9��=!�y�������#��*gM��wϸ?DO
��H�Kɷe剴�q,y���iB�^����*�IW׺���{��W�oc�\��z�-��s����<�;��cwg��^	r� f.���3ܫ�('��=ڞ�vg<W�������Ϊw�s"�D=�sZ3i�IsN�^/xy��3q���2����ɹ�J{�o�F��D\ZN��Cͧtt$�A����G;��]ʯ�śݥ��Lx�3��s�/t�L����*�d0/��8��:.���]�U���bj�q�n�eʩ��tNl�ħ*ؽY)胮�f�H��>z�3w/D������Ja�ilb�0�,�*��e"2ia؆��NiUyS,�+ZvX}ݵ<����;q�.<@��A̞==��{���X��Vnφ��$����횯�/O�Op]�Mvoķ���ݰՈvע��|rm���c�^>�魽��`���۞�Y���"��;v���[�_����������Vx�N>~z{������|��YN-Y��6��<����?<�3�}ƨ�wr��䞍�vI^�.m��t����.��t?2����{yz�h��I��=����<�|�=:=ٻ�׀e�S����_a����*�On=���6Ê�|S��*A����e}_;O{����{o����C�H�o��f▃Tp_�b�6T�6VE�1����v��[b�ꉴ�;{̔N!�w�T]�-���ߋo&�Q]�5a�9���ա�U�A�(�u	j�4tE�����^]���0/g[gS�cl�zǫմ�7��5�܀֋�0�b^sg�W��aL��޻�:�+=f���΀��b�!���G�aopQ�̑?�?X�q=�S�y�ǐp��"5�XV�l�j�R�7V����f���^ݼX��ݗ�,��0C��p�w�w�nN
5^t�7�s��=9�1
C#sf�/}}�gK��p�X������Hc|}���x�/����v�:
�l�ݣ"3m&�1f��O�2�mXJ��\:�{۝�*��c��iCɓ��C�uMQ�� ����wS�*��F�ك0)*��|�=��@�.7��x�����q:<w�y���	������xj��yw.r�^lEN>pm^��n�)��ny:WOx,7.�e�xv�L�� p��������
=ۃ�� z���S��R�m�%Έ�7��ƭĢ�<j�ᇱ�N�;ą�������v����@��j��r��u9��[�y���{I*o�ѯ�L�x��ͫw}y��o�W���jP��c�Bm�U�5m���3�*]��+h]�Zv%�* 0��dl��J��m�u"LMݻ��>�Q����O�N��5�͑��]OO��Q�`B�����PaD?V.܌�
Z�Acډ�w��nhe�G�����=c�?h*@|v��|��spD���x?���u3/��|��^���_�7E��[=S��<C�9,�}�9��|���[5C;�Ҟ\�݋Fnl�z��gsЇ�e��+�mѽQ�,#��z=Սg����0}e��c���j�>����AV����϶zeP�#z�����h�w�k�1��.�.J�����E�Kq+�_��K�b������˴ދ� |nR劥�&!�^VI־��~e����AS���'$3�%=Չ3�.N��5�U\YvY��G�^���A$`=�A���jw�I�FD�ıhN޴&ѥ-VN���4��3� �=S�40�מ�)��K����<�U.]d;h�~�!h�P���lʺ<G��'�^�r��٧J���
p��q��M�n %�51Z�"N�D����Y܉�Q�3��\$�����#���ם{�_���׌��Ӽ�ݳ&���S���Ή�ﴦC���������?�a�`�"R��2G�9�f����k�E�_�hҦI[C�g�8�K�3�d�nv֭�5s��w7�{�;����7ʀ�Q�����.FI��d��~�(�E�v��Ro�ß��3m�������ץ6�{ϟ��eY-9�{\�9������Z��O�]M�{����g��:�A�9ksD��:fHix�M婐�T幤{���)ց��(�}��x�}%�<Y$	3�=^v���ӧĭl�n��ܥ�Zʫ���d�ph�=N�9��x�ze��I5̩�����{���ε�k*	v5ꪭn�����bh�q�t�<;+�w�yaؼG��2k��HڍL��Jw����:�3�DWT{�t�� t�[x{<�\���V�������^xT�˯�����n.k�;:��{��[\��\j�0���=��ط���%ޅf˯A���0)���MD������˪U�H&�:{;�a��	V��c�Dj[�L��V���Cͭ�o&Mk�����R�#j�i�i�\��;����4���Ie��Z����hs��bZ�G�6���v�z��]��a�>�f����y�♨�{��Yv}|�L�ǉ�nvݏn%�
��������;h*wT_�w���{�N�H���)�D	�ټ�l5y�y��Rt������ �0:s��T[���>�Ñ��)��3�Jj�����Q���l=Oyz�n叼�K�=���ITN���h���{���Ⱥ���K���wt�!sۂf��A�z�Y˂���U:�WKK�GGL�I|%�4��+�m��^>>�=�U���8Ox��h%pW�:���}۾�*rOt^�.��9�w��/��ew���ٺ<��B����*�='��{�!yk�tف��rf���@F��I�ݝ�e���_vv0ʔ�����w�����if��h�V�t�td"���C���<Y�����H��N,��|&ń{��	�6�N��GwI�}�=M޳o��)'�剜}�u�0>7t2��Ŧ����^�3w��>��׾SG��_��8/W�o��#8T�nh�w|}��!�k�yæ��U����Z����i�=勋����%)��5�_� ��-l��T�s�ddlN�.�7^d�(~�	�Y��C޴����0g�l"�b{<;��ċG[��	v��|�kR��av��W=�T���<}|:R�	J׀�w��.M�a������؞�>�r5���<����QV@�9�2�\�3!���+c����iK�'�4�C�c�uY��|���z~�����zo���������y�I�&n���9�T�;z���3�'��ѝ�R22�h�3��K;��dj�2Fӗ-d������e�Q�$��X��Ü��(�t��������{�=��8��/7�~�v�^�x��G�>��6]Hz����ky�����w�;��~���ݎ������:��5ϝ��l�]d�led�q�b�V���؃��MD�6UL)j�dS�;W�g=�oL�ػ�G�>"�u�kjw&^ۘUZ\�pM�ؒ���������x�T����7���������mZ����������'E*y�����y_���ju��]�8���/�9�`�����������x��9L��jg5�Z�k�wu�؋&y�EDV�޴�vz;b���.Ä�1���z֢�g"����9���a�a=����IF��Hy ��rN�x�وV�h�)z	�9��:닂[쪁5�����^�aBl��q|����
��Q1��g��z=�A�����9���l�����Rn#㪗#[h'�K��ۢ*z|�y�rc��|}_E�M/�H�:�����v�u��W�h gWszW�b--L��L�]/lF��m!��uz��Mъ5���D39S���4�a'���;�ޙ�R�h#L��F�7��,LM輥xU;�ޓS������%�h���bW��dH�4�hW@{����R���6����r'�N�1LDm�������`8I�WR��z��6Z���k彛���Uo-�cs�����o}^����d���e��r����]����Y&�[�!�!�`�F��B��z�˧�k2yˀ��WYG[x{{����p����3V�����<o�v!��p8�_s��\̄"�+e<�Exe�ck7'f(�38�0��S��8� NJO�h:Nuh�[Z���䪕�Hc-b׻���W+뉴�]«��L��7{��g�>�^ʽ�_���4���X�r�1W���.�ܱ��EDd��sw!�������8ǮG���ycj"�f��&��	L7��o�O���
�.�N�H���bi�'%_js����+7ww�yPoX��!��i�F���:��%]��������c�����7��f�M��yT��}�Z���&�4������:w:�LS
�j6v^�����V\h-1�ӧc��+;r:=��D�9��O�Gn���A9�}C9���Z����vy���\�4�I����ߝn��{���Ղ`��ws]�\�o�QF{��%Yv���~{�׊���{sHC7퍾y�;I������w�U�gsc�(��m�&L�1Ԑ��͹��:"�!���1.N3�X�݃q7����c��ͽ�鋽���Y�{M�Ñ�g��h*ŮZ¿ �{=6��սKw�ă��ں���8��Tt����<+;"��݉5�L�Eƭ)lht�Xt̙̺g4l��,��*�Òv��#%�
(��'�~跣q�z�$|�\�����#�25��ֽ����<����֯m���E٪�wi��V\����E�59�T���	<=y��(����C�^�I�p�;w=�_Y�0�@�@y3��iY旮^4���}�+|o%'�.�h��x�ƙu9�}���;������w:oCw<��%y�ژ����DF��:�����oK�oj\{���6B3�7/�l�84p^��`oe�����&�`j{&�sg�#ch�]�8�������Jo�7�PN䮿I}r��Df��%�Ʒ���̃����)b�����W'���Cw��ù�A��;��9��vBa7��{J���s�5��a�W�78����8<�_������.ku����&3Fo'S}�����ڏ�F�x�{�;��<f�q^��iP�V�9��l�R��\n�N�ǙU�`haL`�a��fqLN����ț��z��c|�������`�Ii�6!;g]ι=�s���>�i���Ȼm4���ު:�Y���wZCd�%���`�f�_��@�d���^��;v-�=��{%��7b�>���k.������z� <S�٪�8�,G�{V'���x���ȳ�K��j4#�;��6+��iF`�$�i��4`M�b6�zhl�������܂�e{�D�c"V����j�o�魎׸{�D:�1�4&��G��t��-P��j`��x-WQ@
v�h$�\���n{�Ġ��U�tz�Ћ�h-�)��;���t1�l�~�n��51��U�OA7���͈yd��g�`+=u#Ν����3�ٗ�k�w�r�ӵ%��+��N˛�t��}(�?)ȏ,j���/���S�L-�����d٭e..�x�;]����Aۊj�}{&����:�˻Q"[M�-��D5-�VN��s�m�����rZW����+��<=7����M�x	}�r�O�g���׾�uY���K���7���dU,\�.ˌ�9�ǚӮ7U�gm��H	�*����R_����o{���x{��(��=�� �ƛ�bzN:��I|+�yj	��1���{vI�q�_�S�Mn�}5v�ދ��4n��1�ԇz�M��PWG����}��-�ov��>��_�";�iP(ϳ[6��bw+#o::-��+qQh=�	��y�6�N��X1�A�:�ϘѸ�Y��W�.�5d���,Xoڧ�C����8��©����ڄ�8�r���0��d��ɖ]
��f�u�/JrP �6��*7�}��`�vh��1��6c��2v=�k��Ǻ�/\%s�}�A���r#BTa��mh��)���x�m��[�99�;��`�䷱o���]<����.J �8vO-�O[��Ӳ�Ǐ&����9r�#B�M�īo�n��+�RǣR��L�� �{GH�NH�����x�R��P�,h�(��zTV��-�{��6'R�2��Ox�[�^P�3ύr���[�簟X#�[����Y��=)�q5��B�$��{�ė�x-�Q����i��;�S��.�����o��N��ZW��������c�4$i��Dovk~y�zf��C6 �i�.�7_��ǌ�>/�#|f@Q��f�'��s.y�f�$ ��ú'L�$qڂ�J}"<zF<�~����ݜx�L���f^�dm9T�����Ef�D����Ö��N�Z$X�ё����ͱ7=�:���.v���;A4YwZ`�\���_o�%x70x�����{O.�@��{�L�`N볷�8��'὾���"6�U�g=ɷa���֙�Ѣϲ����=�0�@�J+��� � "�ПB���<��ub�&=Y���![�E����qYr^��yp'%�V�ٍ��ܕ�ø��M���A�=wKc��7��K����Gv��kF@D��^փ�����7���B��Macycq:I�����YXܲ�F�	�Ǳ�I�[��V>>�\"����$ ���WcSn{$Ŷ�p�}=۱ko]�}o�u	���Z�{�!qv9<>}^�Or�ށs�N�˟n�r�}7���)R�-�/���~�>�ܯs��������of��n\�s㛟�s��r�=�G���6-ɰ�9��]/x:���/!� ��»q��F�a��n�l[��5Sm��vu^�vm�sN�u G<n�L>wc����v���/X]�{<��[�ٱ�9�`��1��{M��H��=cQ���OZ'$�[)�ro<�[s���Mn�J	�n=[�m���/Y�tD:L���B�qd��b�a{��^qb�a��.�;����[.�m]�9�@����u�)ێ�Ꞟ�ݰd^6�&�T�=�������Ѷy�\����\upy�y�y�Z�m��=�8^�x�wL�svH� �눪8�E֌��M۔�:�����h��:�u�cٛ��˷%u�ݸ��m�aϣ<�Z�]=�t�>I��a��._m]�mcI�l�[l])�S��=�G#�.�ۮ,m�V\�k;<c8�<q�E�����:��ㅱԥr{]�ju;�[���E��vN$�q	�b��{&3��:�f͢x̀�)}��q�ݽ�,0�m���ܘ���۬�k�s�6��qN�7*Z]�ݎ�;u�s˲h�]7��ۮK�wa�n��]Y�s��h�Ͷ�3�U��9�۴jؓ��<s��w �^Gh���!���U��n�q�C\a�q�y���P�=��8�qx��Nݦ����{'c���{�8T�˽.�a��v5�m�e�k �J �h�HF���>�i븸����:`u��YT�!�6�CC*������k�҄
����%��������z���*ql�ݲ��ܡ�{k��͵<�wn����yz�ZsS�米>��7g���d�^���dwi�E6�&�7&�˕b���b��c��S�cЏn���Y`�U�K�Of덊W�qrv7OnDq��FnG�\Y�*�^�p��K���ӽ�$��sÓ#�.��;Z��T:5v;z��خֶOj�K��&ˣ��ܹ�P��v�Иz˭����2u�^�p��M�η̭ٻb;z�4W�9�6�ݵ�b���wV�9�۶�NL 839�J.���n��K�����Ǌ	��I�o��x\t�	�,��U���o4��)fKIh����mS��WF13�B�� j#�A�
{7X����b�XnM��d�(�CT1T	{� �Ν��D�4г<8�w��D	��	3�O7�=�Ll��ӎ�fxl��WC��H���5������O��YA	:�h~\�ME��ͣ��E��9���4֯�:�$\9ܚg�wt��3w:Z3�������[�H�@f���p�&y�ͻ�Bma�Sz�:3�L�<F���{���}�,��]�D3���n+�2��ݺ�&	�^��׈�9��z�i+�|I����f���w���ss���ݵtȌA=2/q�>'p��o��<�hEM�پ{�i\N�Z�܉6�&mÔ�8�4�&$ǥ�]��r���g�J�����v4�����S�6��Tѥ�ft��Ǉ��/���9���p�O�soc{�ZG�n@0�/K�'�N��zS��/�{���y��w7x�
6��U�E��J���A��}΂M�N����t�(ˉ.��Z�WDm�XI�Dԉ���xf�A���#r
z��w/^��I�Ӳ֎zl�S�6��� ����,�J��&��ƔL?�P�:�^[�ޒX�L��$B�r�s�$��-��=}�����a���;����d��G�)w>`S �=���ٜv�3�y�,�V!K�N�1�3������ٞ���
㓃��x�����=��5�P���ݎUKh��2�����X�FM��$�����sͲ���9�Ūxw��'�;;����N/tݙ���k��)܊�I�cvU�*���v�'.�S�1��e#�-Z�> y��Ч�2�=Fg�ֻ�w��K�it�M�)���b�ݝ���4[�X�!z��=N�3����n����������8��]���/ؿ`��mK5�-��y��=�j����p1�s���G�kя��t{o��Z�8��:��Ͼ� ������M�x��K��9z g��I�����{���K�Q�J�'=��.��������/��ǽ�O;�q8�89�EB%B��ezfT����]F���{�󧧡ì��v��wI���}���rD��B)xĤb&KN��h8��Rî��#��ai��vul�$�S�"�F�V���Z_7�k��~�8sjzv��Ke��x�#�}6Zt��IqE`�N���M��u�|���U����ѱ������wy�("��)`K��^��9#;�N�x�pc�+�>��YN�\��V5R#U]�KӃ��^��a�8q������#���\9+5t�	k��M0����c�o'�	����⯡T<���}5����75}D���iQ[�&��l��wmЃ���ݾ��W���������p�O��m��#t��U����vI�G�̺~��ϊ�~��X>Ir���y�R�7���1�;�a4S�f�.�i�Jl:�q-��h�
iPbO@BRb���륺�[KV����^}�|���\;��q������" �&IL���=�� ��z�\���������F�{c��ue1�A�$ą"%�dj�8ݝ�����N�Yճ��[}����ѓ"H�R��'�N�Ꮍ<���[[�e�F��8���#�f�Q���>�#�t�A\D(>��s�����խp��O�8��U(�D$��3#kk#]������=�'�rz\���V�Êp��d����((%$"L�)��յѴƭ��������vZ*k������~�:/!y���#�)j�ܨgw/^9��#v�ÇzjN����姟:u��3F�w�������qdld�<����Q���e��$�&ܡ���E�a���<K�{&�(��s�Y_����Ӱ���'�H}P��<���="��;�������9o��IkM0�}�J-/��:uΝ&��S��� =S�=�шl�4Z�Il�A7w��=��R�Io�bt�"_[Ef���� &���!D+�s�7��v�p����:[f��\X6=�{un��n#zօKS��Ӻ����s�Ý\��Lj�/i���.�����ؑ�!@JQ��g��D�ղ����=�u�i�k��;M���� ��w	 �
�����-��5m��;�Y#�3�v'Ns�pu��p�' ����!L�[����ģ]ˡ���6\m0��p��ֹ�_6�YUO��̟Cȑ2b������P$���5��iۙ�{��]��v�T�F��wo��&�\ⶩ���q(��q�W~uw����*|�#&��dE��{VkC���Xtϙo&�;�rX(ea���}�{����<���R u�(J^f�yŻ��Z޵���˲��մ��C����'�t@Q!$�����r^�S�A�M2.��B�� Z�ݗ�V�K 9����B�X�uڈӌ�����V���[nSg�� -k���kw�	]�N�.������t�����_.�'�X��q���P�n�E������122\�޸s��i��{���}R��s��m6�R�%#"0DB�R����/�nC���.66ֲ�5oyi/ۜ�әϺlru�����2�y�6��[|=��:i��s�Sv6��ccgq���� �Ś7�|g'�����F�ڻǵ�Y�Q!Q�Rb��u�&�P�z�#Q��ٺ�ø{,�mr��Z_1�N�9���nۻ�h;�0.S�6�丹�ս�pb랲[`�n������]q��wy��nWcu2iTs6���gۚ�dW�����s|k/��p[q�۫��&��&�˻�˱s�v����r�Ѱ���j�Չ�#�������d�o���X�X���v�~w}�>\��ry40�]+�v`ޥ<ֺ���x枺N���v�A�8շgG]�ҝ���v���A�&��%���OC�p,<����
m�<�a�w�|s�x�G���{��n0*�����LD�0�en�ˮ���;�?vx�4wZzS ��:�+�\h:C���]�����tdK ��G?>m�0%L�N_T�����kkZw?����n�z];�4(�	�$�$A2��Oe���^>�s�Ѯέ�����G���æ�� ��V@���s?o��y����� �yٝ|y:�q����PR���O�J&F�������|rs����뺗[��x>��i�uC�
fLB		��ʙ���+u�[]���\��:���s���ٳ�.s�Ⲩ埄YZ��V�.Μ�vx6�'��p\��l�yjQ8�c���@0)�c(�#j/^/����y;N�[�k� �#Ë���kk�Ph�^JbbJ���2��OXuo��A+�KL�F����E\ka
���A{�i�h	&LR�å���d3'��臹�WZ�j�0QA���~�'n ��EIF�e����A��� �>���Ĳ�26~Mq��=;����7���Bn�ᜊ�\q.�@�P�^����s���Q����u;[[�w�<��>"ɓ� $��P�13=.�zXu�V�]�7�<5�C��o]C��k���2�̘^Q2�Llo^��.�W3�����������}�~��s��jEGdR+$��wY���[]�(i����s�놭��7;[:�uv=u�T�Kj�Y>N���L�cv)9��ڳ��n+�f��.۞-ǽꍹyݙ��s;�߮��әż������{ݏ
���'y(�!D�Ɉ���\�9�cxx =.��X���q�������3��j��Q�ʀ�
aӒ�x��ؖ�p�F�$k��fd溞��͌�i�D�9��U>�4�[{������Q�n��	ws�/�[�8s��#2<�<:!���ِ�l�����hvl�S��	��_kiG�{�������1�u��8IyP{���x�S�S9��}a��q�}�����gr��\�g���Q��Ql�u�U��ޛ�N�mt��d�a��������p�b]�㒦�)U�9w��9����iM/u>���a�-��峱��{�lD@�1�Y�uٻ/����-��qΉx�f���;�L&妩��������&�i�$�+(�������+uƭ���=��'�Ϻ��unl����&�b��e���.qo�$��t[�N\�o\���R���y�Q�G�>R�(AQ2]:\�C[e�q���~��y:Ll����F1I�B$A^^P�����{���:u��˭��������5��/�H2{�9���z�����������=��s�ѐ2�C������вk�1���I�<xI]�KU�=���O>�3�}眤#$pC�����1�C�iƼ1b$�Q�D��|(h�L��$�5�1����hGY���I$#��3�<��OE�	[�r4B)$��6sw�=�:��\k��B������;;]�������.}�]�S$n7m��I���E�'&�V�l��'���m�UMh%nJX�����s���F����kl��;�<Et>���H؞��[�Ԩ��ٿ�q��G'_eC�[ʜ�l���x{G��K�1H�2fA)����}�8�z�����x{��<�߬]:k�1�xx%��M��{���Փ��C�i�P���$kKg{����Ω���29J���f���xO�:c��9ֺ���FӇ[O*Q���7[����93{!U��8kc�bц^Jbo#�:r���� ���j�"��1�Oi46:�"�	j�9x�L�%�RD� �M�����������Nw���yx֢ޣ��X�X� �G��V��Nv�h�b�gu�rm�N��ݽ�L�봝8��ؿf�J'�럜&ٜTm����Tk�ٕ�zu��ra\���;j=s�4*�I�<�F5Ί��)c5Brl$�=�Ω���6-�����.����R�����9���n��<��kckɤ��Q��۬�-���1�,��D�T$I�]�r�-��he`�B�(�@ �3H�u!�����ŻGj�,����7�Ya���	\��ۛ�ɼ��](�ꪕ�j���������^I;�+��[�ػN"A�n�3��������Z���EI���޾M��w��m�:?�	�x�S����LL�
D�)��u����{�=� c��8e9+w�V�m�>�����!AS�IL�[<��s��L���=���=q���gM& ̡1��:���xWMw�;ɝ���,9���}�Y�|g޺�wT,*) �͟�ϲs7�ִ����u������\j��s�1�ff����f�vn�>��;��:;z�Z�e��)n^��e(��=i8�d��N����[/S��eh�K�OOqp綼�b��!��-)y����Ns3�����M��"+Qma��.�������7Ӝ��(5���s��}Ou.�u��!��d8��꧴�VgH���1���=Šp*��˝���=5Z.�S�gSъM�;�d,�o�f��<����FS19�qg�j@V󺌂x������{^�|2�)�E�jϜ&�>��S�/jX�����2��ʃ12�#2�JK�Y�Զ��5�mw��p��?v�W3f��g>lR���I�����gGe��G��ll��{��l���x/�$bƃii&���yz��<<7�t����Z�����e��	}P91�z�@7#f��XXP1ۣ��rޙ{;����C]:��U��MBfK���d9�<놭���:�z������i��:���eB��h���o���@d{�w]N��Z��mͧ�zE;lt�[
��I)	R�]�����mKN�x�~�9��D���W��n����~�urFݷ7٬أ������RҲY�PQ�#��ݢ\8҅C͍�	(���;ؖ�PutC�ٿ�{�|���(�-|�nt��zӑ�����w��OKϚ��xy�sP�0{��p�&��Ly黾y�Rǀ�M���7�#�dj�|��F��`��Ơ��N�9��ip�˨�ݻ)֭����]}oC]�
/agtF�d�Ņ����7�"��7v��y��w��״������������Y�������2[$\�c)e��V�%;0H�S&�K���b��P8�T�$��mY��Ӽ*-ꑀ�;�5�Y�<g�6�U���r���z�C��#��~�����Q�"UZ�H��v)o��t��n�3��KdC}� w'��>]?7�wljǂ��
�O�[o�'�1u9�6b��I�w����N�4�pWK��N��Ǣ��}z�Gh��R4������M�{U]��7ks+�T�Z/��a�4g G�[���	���՝C#/S4�����W��S�n��س�\�DG>�7�b	����v�.ٜ}�x�������דۂ����G�s��k�&���k2n��peudo����r_";|͹v�뿢�9b�YNo�����D1��+�GF_j>��ܑ�vu񩱭4�^�7B`��q4^u�`��=�����q�3N��s�7w��#��V���C��R�ۢ�6��)r#j�1�����V���܍����i�������a���L�Љ������ۮդ����Ǽ��AѲ�C����Kp<[q���4dbђY���y�����eL�{�Tf������|�@�A�NqҌ��Y9Y%�͗��'^�'F�3���6OFd��t��y_G.B��'dM%,W}���PU�x�sͩ�4�J�kx�~t��w"�M2ɽn6gJn^��!�ݼs�G�=�ۛ�#�T����;˳{kD�n��Ooijn�P�$����zwz��7V��o=�nA��7'�����_*�˥�=S/cL�e���SLa�+jf�<jQ��}��y�{�_;�^�P�M��������2򄹍vk���M�8q(#�sʮ���%�Ã9z�k��c8���}���]�6�r�<ո1�2���w��/�s��%M����b��L���dl�&m7,\�MF��c�N����1�M�11>�6�w$��r��N}�4��x`h��v�f��\v�����Cb]�ŅEV�<H`�Z�>���^95�/և���zgu���܃&]n��q����{[h�t�6���/����{��OoH�[��ˌ�Mn�����}� �{�x��um5�;�Y�ƽ-�w"�M��0VM�yDSD,ۢl���,4���=��z��0sCs	t�x���)u+g�^�`��d��8��ׂMxs���A��P��_3���&��^�s��-nu���]'p�{�~�I���띳{��cth��՛�;��Һ��4	>��.3�{��q�_t��o`V�ף{���={��a������ބ�Y���B�H�{W�xG��=#@ˉBx�駥	���Ëte��d�@�)��)$��&�3|lV�I%�ҭq�XͧŊ�RRU%3IZv��xN�ʝu<w�����/=��uʒl(d�
ě�{qI62e�3)fgI/���3-52T.�q�ŻD������"�i�J�5	��m�ebK�f�J4��E$��2��J{���+���v���y����D퓦퓦�)aީm�Y]nƯ�#��e�R6�<��j�q��`-V�UD*7-���*�K��,�(�D��/I3�M�MF�5�;��V�BM��2��Ғl	�	6F��.L�'U�t���<u��âx���u�y���������TV���P��&��N��9G�W}�S�/.�7J��]�\^9v���]�=.غo>��yr�]���q/,�2�wyAi�	D�u*�4���Mf�����M6���P����i&ҎI:d�-�I�{��n fKD��9���]kIWƒ���d�߂9��f��ӗG|:n�%����ǎ�|�x��|�i�]�Iae��M1��36����b1V��
�{p��u�H�$i��ӗQ[�8���c��"+{%ʢj:�Y���ے]C�NqU�u��H�V���7ߑ	���>ӕaZ��Oϑ�y���0�4M�!5�b�}έ�N��.�Jî���cgv�����i�%S�ՂnIO��Re�IY�eB�mb��C�'�^�OD��,��3�n��2��vG�r�<�s��q�}�����ReℓH�fY)��Txd��d�>}��v�ޮ�D<r��{��=������qj2	�)/��\YF�c��@��̚����h�X��[�h��%���#7�}!�t��t��۟.}<Q֜/�;��{��\3@�d����J�	2T�4��2�J�g�ߊ[ɛZ��@���K��褛�-	)�Ê�۞Wl[�.���G|�R�n�W���dp�@�ŪS.k�%��IX̺�T��h�`�$�+t�e��c$��I�:��d�kh���o�2mX���=r�k�,ꍀ+*ĕ.d�4�aɛ�L��6og�����K'�on��:jv�tv�ۿ�>��髶�N���w��.Vh�Q�j�� P�"\SL�4��4��3���Z&R3aG3[`�%Q݅&�K�M�=�S%����Q�;�P���@���#�������}y�q�+\��zGM{�Ei���Yq}Z��h�rُW@D
<�2V�'��p�5�&BWl�JJ�p��vB�$|xd�����_��{���H���G�bх�[���Y5�i;Eúm�m���pve����Zf�g\F���Hlv�ڇ
����m��n�n9u��ϕ/-�g�Y۳{az��Dk@�J������N��5�)2��=s;Ƕ��nۥ��ta^�����n��ƻ$d5]���݅����}$��.ݷ�l���v�����s�c+����^6����=�vs=@\O�
���d��o���c��	�3���q��b��_w��Z��W,(�������^�m(�0�@8}#�n�I��-���@�aф7�/;�:��S}����t$��f#J���2n��#��c���K0i�U
�V��i,�d��4�37�f���$�e����t�KmuÎ�;wt�G�q;�w����s�yn������,~���:7,�KEni1��%f	X����V�3S%�	h���\S7�bm>z+8��V2��������_������ץ����^Ru
MOJ�eF�*'��zє��X�>n��h����Ж�$�7�雊xf������^���K�rc��-M I%��Қ��H�̒�hd�I<��(i�����-,Kn���6���̝7�����4�Fk;G>&aI�"i*�����A�/��u����3ab�d�3;6wO�����EBd���L�P��5��4ͣI�VrIFwD/<;���E��.�SMv�1�<��Nc<n�m�"����#�JcXT��aa")�-M�4�3X�nO}5���By�פ�@�3>n�əٕ�ch�|?w|��m��ǭcS|ן�vX܀�'.eΟ
,�dC�4�r����|6څ��U�n�&_EX��5�I����2��̪�e��0�3��3ē��T�vgQ7��i�>�"6��3��������['�g;
L��9}��v�xҞ���- P��'L��\��=|���E��M̜e��7�*K"m>ٿ]H��İJśu�L��e*	�7�R'���q��'�����)�Xݪob�	�M�	nMꤖrmd��X͝�礴�������=3`����o����@� V���ɝi|����R(��f~���(�2��L��,��su�$��IjgoފK��њ��J!����"zJb*���&�e���+Fk�W$��(Jwy𦲄�P����Ih�Ko�F^�3`����{KY��~�89
U%V*�`$�E{[���f�nn�m#��8�L�-���[��\�(0��}�f�<ү�%�K��<g�2��S�O�%�@���+t�LؚE��J�����6�h�f)8t���	��4�U=`ʆ�V�9�T�v�KHz��q"ZX���IiB�5����e��P�K��}p�S$�gr�榞�II�P��ߊZ*�� ��Mq��蟄�Ц��[b���ejپ��G�yҤF`PF}FG�'"�i�A�{��Sf'�O�[�(����Ƀ����H�C�{��mk�vd�[(vq��dܻp��.���R�m�ZÉ�k����t����<�xN���ڕ����p��g�g�I��)|P��s+U2�4�/����"�T�R&���Pg2X�	`��{��-�-ί��acaCf�{�4sP̱����礼Aᕍ;.�TpIA����*����,�Q F��2���I�%cJj͞zn	|X��z�- K�Y{4�J��M�}������u�d�W<�Խr��Ó���y;:9�;v�u���P{K���I�n�b�2�=p�E�+��襣Hͅٿ\Sib�����ɕ3;iCh�����xj^�8q�׺��#�b2�,�H|�Y��T-�o�hk��[ޚe�EB^ί��K`�d�E&�rM�%�ֿ<��n�#�H���ǋ�|zV7�k�X�C?�~zl���$-,O�\�¡/	Y=�t�h�L>�=.�FV��!�Yǯ����RQ~z;}�\4����E6�L(L���RZP���^k��N`��7O�ם��P�U`���@ܑ;���ί�GߡC"��A�tF1N��ʯt��ې4���lZkޜ�<�rhnT�	(���q�������������M����=�kh ������������W)�74��rN�9�J�:A�D�r���c}�5��������G-��ht��%&<�P�eC)��U�Pa��3�	CoOz�m$ZP�z�)a`����k��+���U����z����b,o%7�ŷ�!��1'o(C���U�Z�㧵;Onu#e��.��ֱ��.4��?�^��ޒ�ł���z������h�7�LK�c�K���n|����f��d�|%��׭�̜P��o���)qcib|��)-��P���M�$��O�=|�<�����2fa�j��P��8���1�ҴS���J4ql_t�n m�s���łj�քj�@�D�<�Ma�I�%��WzkD�-(O;�����^��ޖ�a�5�:o���zK�P�Q�RxQ��*�f��D��Y�n�Kh�l,��'R��V�%�X�[�L��`�>n��i0TȻ���_��?������{:���ݭFxFv!�/�k�p��̃y��=x,uN�P�#�>�Y�y��͎!�V�H��5c��5S;�vѷ�9��Y띘��ݭ���w9�E��;��F��8y�tD�V�9��R��ɢ�v7룶�\��v�:z�7&lr[����d�]a������S=@u!n{rv���t9�Ca\��uB�$m<�����k��VV� ��c%u94&�5���tׂ䇬�}ͧ�nѪ �nz�[	vF<s@������"��=�(��.��66�D�lҹ�:r�A�[�H��&��r6�{~��/wZLM�� �J�a�&$pax����-�����Q��|�}�۞����\�q�����.
�1��@9$��]k浍.\�Mi"�X��[��҄�P����[6	G
�"�������ԗ0R��ӈ��� ����u�ZrM�'����utSh�6���M���on��KNfT��4f���9�B� �K�f�EM=xjEbe�։�XY���Զ�rf�3�����KKh�<�s։H�Vds���mP���\���奉.=���Ō�X�Ϸ�l$Kc?�O�҆Xs4�=�9ܩ�e&��b�S0Kĺ�RK��UT�F���n�kF��|����-��t֐%��>�~)`�X/�nw�Z��X״�)��B��BJI8�u\'hq�b�gcA����qy�0�;���]�=������5%�Z�[�3�_>��w�{����rw�
��m�ɗ�ƅ�������׊4J��+d&!L�BT�����>�����M'�+���f/�w�H��W�7���U:-�4]��՝!\[�[)�j�j�͗��t�gY�M=�#�g�04R�j6uVU_H�9�nGN]�i)C�7�=�|q�c��y4��; M{JXˣj��Q�5f���I�>�(��tPf��|��Mq��k�%��iE������q�>�R�+Z��IUFV>WmH�PabY�[4���:d�E���WM6�-���қ���gz�DM
Jx���kI�(�5��[�-��}qX+��e���X�rM�$����(\Y��r�G�$'���䩑�Ua"��O�����fmIB;���p�KK3����ł�n��R�C�X���V>vy�����MTF+x8s�,��s�E���ۜ��^� ݮ7����}�I����3��K�cP�T)�U�����ݺ�������\�	-���뮚^j�־|�}O?2j�R������K9�V�%��gw��qf��ί��V,(�e���5%����u�	��^D�ʊT�5@��O��Wj�,�"%�E�������O��̻�=��9j�="�ͮ����]�=�/a�I�a�D��-��IN"�$۵3[dr�u�Ds��b�#�m��+�<Cy��ӹȩ����丝 �p�&��^ޘ�h̅�(�]�v���<����}�x��W��¡�T?��RP�qk?�'�\$y���j+H0�f��u������U��aB�ݺ���L��!>��\�_5֗��H�"�q���30���#n4���aG2V�<���K�>���[֖,��_M`�,(�M��~��O�S�9慞�-�Bv�ɭ�"N{��=��;���Z���[�v�K���w��I��6T�P,,��?�~z҆�P�z��7���<-(���ip�h���оR�E*��JJ,\x��5��߮w�2E/�q�¯
F��7▊L[[T,93y�Th�S��s��Q�)�%V�-��u�Z(2��ޛ<�K4-<=���i"^���[֖`�b��"��A#����	X��iM���j4�q�} ��
��b����߹�+������Buzئ�"C�,b ��'�]ǿ-��aF$>n�+�����V�T��p��s��5G�}xG%P�h��֦��Hl��|�nȩ(����ܑ����q<��{w���V�|�8��X�	�������zK2kۏ&�Y��~߾��q��̽����!`8�
\]|'�ުX*0TrM4-�ޚ�E��S�*�H�_��U��9$������r��/�[��+��m�k#b���}����X�]�{;=,��v��om&������4�uv��6
�ۭ����S��rL铭�O�}��b��E�xR�C��z�z�Y���{qXs'���ݳ�)h�XPٝ��0�z+uV��P1-ƴk���܅<�*�fi��gm}4�TaBmꥅ�-d����\W-���ΫB���d\�,�#�Q�(���־֨-�徭Ě|3�g*���v�b��q�IwZ[��=�������R��$�
�����5��߭�Eb�_&_4n�zj�b����ްV,,�yߢE��*"�4C�.��0�?�>D�w�԰��wEWZ3��u�*�ܓ��T3Q�8��+/��������������q�$J������\�}tР�����o��E=�T�u��1��١c���Hw]��Q �	�g��e�`k����vt��M�{���m�����V�*�om`�&��ks̺Ss��$�������v/>�E��ú�d�e^� N�n�Z���>0�ec��g���������"˟�y��l���M�c�<�Sϡ����fy r�_?d�7I9�۸P⭚�߸g������X�K+їM�m[��)]�	�u 6��Y�q�/�ٴ�w>,B�~��{� �L�9p4�(�Y�u�o,�=E+��ز?!�YG�������%F�I�	����cɇD����a{fp���G9*�7ܖ�F�s����l�Ԣ��{��˂�e#]wD����D�n�6�(5=��Tq���#�g�-��pkY�)b�]Jj����]��u���6o���R��)�r���Wb9i��Z�����Iq���M�ȸ�#�u4}2�>]��]����Z���;��;���+Ut�=Z��Z�S7a1��iܚF���e�{)���?/���k��Zz^��o���k�����Uppګ(���ޘ��Ǻ�YD�X@�F�G3���Y��� �<�Y���+�=��F�MC��^�S-GB�y�A��mY��@/�v:�����B���8*ӓm�\v���8k&Z�	��"��*̤ۋ�sû�O2���\c�Q��]���6:�i����S�:j'fK�vޘ"��$�^���@����BzΞ���������s�����v�ks��Ե4-۶w�۟k&.��v�`|]sbY��S�]��m�R�zl]�-�nN��M��ƚ{�M��:�q۬���u���Q캊�]v�B!��ˉ��vԁl��l��n�N�dwS�i�)�hn�۰E�:�����u��)ۭ�v�ڸ����Nz0��@QN\�	<�V���r�wm��bR�	5�h�i�#��ˑ�b
�dCq��Vb�t��Y�<��	��kl��6��s�����<f��Lr�Vu�ł㪄8t��8�>y���h�v�]���)��nL���c��w\��7;$��=\��ƹ8�����v멜�@ݴ79��r��[G��{G�ݦgc��&�k^P�^<��z�y�a�!]�ɇI�vrֻ�_[����<i���OE;�f{	x7Z�+=�P��Θ�B�np�u`���vN�E��\{<�흺]\��3��]vT�9�I�s��;%��m�M�0u�w%|?}�n����Gɜ(Ix�X��{j-S��nm�r/rnhxv��1&�`��m��������.Uc�W
\]�7:e����=.�ͱ��㔭���b��l�M��V���p�rʒ:�Óym����w�����X�jTN�s�8|�[�i�Ѡ�D)�Opǭv�F���]v���/]���Ƴ��c6W>����c8��)�����b��a�y��sT'k�x�+�yܽ���%��Ԗ�����ˉ�n:�8ylqΣ���W�J����1�K��:� n���t���=F�ؗ�.�s�����)8��М�Ò�ˎT;Wm��2>��:�g��ABm�容�p헆�qǷO�*zy.x�� lw���x8�4 d7���*댬lrupu�vwqt�6M��fe��h��Q�6���[V�Q{>��9!��k���Ǟ����8ۈ��gw6�qfBuٶ=���\aNxgc��`�YMѻc8z3�q�[[#]��G�[�!��nX9�Q��dMi��A'��0nN���r��d�Q��E#Mr�����m�Ņ��I��;S}گU|�emw9=Ξj�z{���8S����8����ٽ�.HH����m�u�{�{W�???	P{�<\��=u�Z6O{9ׄ]���%�����-��Q	^�kk^]�2�P�+M8;b]�%��k���pn��յ�U�u�l(����ֈI�wNB�]P.'`�<�;G�f2�c3���n�G.���d�����}`��,�|�m�}�{H<0��p�[�X���"a�[����q��Uz��a5{zj��=axC��y��bE���r�4H�����둥�=����'�|�Fw�v魯�n�>�;Zb��`Ȏok���.Ĺ2h����GHa�v�y�f���S�!=��kԽ��~�^E����M�`~�|7���o��x�A�>ˣOh�af�ۤߞ�:�����.���jK:�nY�b��m�ժ��nv��o5�ͨ`ڮ:7��jx	�����|7����<\�ny|d ���4��m����T��������6%�`�u�$Q�&�g
�A�5jȝC̬\�[<P.ם�����fܾ�����h1��	���{Ƈ�q��h�>�N5�鐬�k	�EY59���Moڪִ���|znz�/'�����{�'g�j������Q��p���6	���M��1�a�2)��U�Ӡu`��K�5�xW4x���]�:�c81�m�5͇�J���~���#A����<Y�g�.ս<!�Uߖ�=�,\<��g�OnT緮��z8ӎ�����	044()%E�C���An�gK�Ccm�88�8��ՍkC���۱�.��uٹl5�`	{{�uvW���f��by۹��4����X���nu�Z�� �ǩ���=[� Z� +PV�4��y�fa�ܚ��񻘞p��v����r��l������&���w��1��FV�N1*
�7�Z��n��J�'��ig���`�1�OGg�r��.'���`X��dmV���RW��'���������X;,FV�~ȫK7;ی��Q���D�+nX:�z�*ꋆEӸ��ܧ�$�}��X��v�Suc%��<L�p�\+6+x�����ih����_�62}>	X�f�ip��Y���C� <K�2�T,,O�z��3*L�F�>��R. ҆�u�,X*=������i��j�D�.D�`S3T�!8~�T�F�e�ag&J�M/]��ZY�����P��j�˺"Xx�5RI3�lJ޷� Z+=�R�Ņ����Ra�5%���Rҏ
��sގD@�	��DL֊���uZ*ɕ$�OwS��I�]]T- ��>�j�G$˭�(� !����" �E��y�\��u�����C��XJ�jX&2�m�sk�`�����r�YB����u��~'�L]hxQ��e,$�X����s&�m�������ZE��Q߇`�$D�$(�
&���L�0Ti{ �����*{��nk�Z�Dެɸv|�2���k}��_Y`ȫ9A��v�qd�_F���F�H��q7u��š�g�@�U�s��p�����y*���9\����ӆH��3��c��wEݤ�,	bD�'�w(7s���u��8S|Ԟ7��������}��1�}�ȭ$X*+6+I>n��\ͪ����������QP�Ŷ>	X�&�kK0V?���-��2}>{�+�&�nw�T-,���Z��	�95SX@��f�g�Oox�$m(��})h���O�m�aF�';�oZ/�^�{ï�RHӪ���3�c\ۿ[֍frN$�����46�ibm��҅���7^��ag&J;~�h�9�]^��曠�]����g�V�Xù��gN�l��뉸G�ܦ8�b�鍹�m�;�5X��ʖ,��/b��`�O��j�$�6���Ep�ҏd�(S1�����if�Z�93|�7�Gw��ť
c�iKE9����Ik/�k�Y��U[���Q��`L�X����\E����4ȧ�deK�;Qi�k�����v�9�j8c7$>�_sF(�����Q܅�r9��q�b�ZA�o�n�'���u� �fb����Lx�:[�j��'��%���iͿ�SJe=�f����Mvz�U��� �����]�2�B{��m�>D�	�Þ#}�д�bn���F������a	��:�\�Z�}��\)4��]ʖ�`�Y��5��c.L�4a[�6)�?چ�����K̕��I�̙x�Y�ɝfǾ�\P�V'�zX@�Tln�ꖊL(䕛������:�h}:8r�]�ʓv�vκ��\��j�;W93�vD6�c/�Ѧ��	�r�1H�-i'±w_\V�`��N���aG�~��L���_I�m�д�K�-g�dr��EP�3��ƿ>���~IoYV�<�z)h�҇�v�m$�X�/nii䐗�׭�~�K=�R��v�"͵��̊��A���{R-(�o$�Og�s\X�Vz;�+<��& �""JZ)3�52Qe�o���/�����(�Q���+Eb�)��FWd�z�n5`��R���'\YK�GFI�+�r���� Ω�O�F�+-���Uw7x
�D�1 OgX��CP�r+����!3G�n5��wb`iћi���='ο"�� n���ϹS�bqP�<�\����FL��۳L�K綾s��)ڨ�4��03\x��O�{�\�R�T���ċK��E-�P���KJ0V.I,ߗ7Ĺ.�m��Ȉ�N�ыh��v���k���P�sT��En���"u_��^e�R��](�J\��־6��h�XX���Z(0�fm}Ts7��i�0W]��/-�u�#Ht!�T�R�T���Fm�k�Ó(e�O��祤�/��߭�K
��m�aəٜ,Zx�� ��1*H%LHV��(�/�hZX��oF^�ag33�Ѣ����$m>=�_E6��(ݴ�F��wyB2���>{I=(�5ޞٞk�ֱ���:�(l,|�حs&�I�~���ϯ�^�fEj�+42�8@3��ƾ~ݯ���a\�Z�O}�ԴPiC�o8�dYݗ��"�f�v�U�]W[�p��֟��yo����تVzhr&D6IQ]��c"t^NcCH�wڬdn;��YA�n��'�S$�4uG�;��N|�j�����"A�(To9)u0��]��FsE.kS��䆜�mֵ��{6��Z���Ϊu��í�j�j4��n���3r�;l���oku���A>�6�\�l�	�.��ɋ�)v<�ȢO�cK�;=;�uۊ�:*�a��e�㈮��`Jأ7p'k�TDr{�[�n$���M۶���7ϋm[��XEՉH�b�c�x9���b�~���������>��+���ru���͚ �ϟQ�ǆu_VV�d�$~�g�7�ђ�s���Xo'���;`s�8��i�K��I�(����p��; �Qv�n�t��U��q�"�1a��Aa
 �4G��'&b����¡�{�P��{ ��
�f�~&R����x����1����v��e�*hv��Z�ܽT����X�V�tWh��|�T6n��V��jeQ���'�9��JVV�	Lƺ���z�{:g]k�~{�ߊ��d�2u����Ωh�҇��zZIdYɎK����L�
b��,��+L�����ZQ����h�V�Ҍ9�bq/:�߹���lD�Ä�!L#̽ib��Nf�R�Q��&J��V��-$�T)ͮz��oЫEBIQ=����N��	C���'������`� 
1DR��P��`����z�0��m�7%�s�!���{�f5�$3�:d���Wv� 4=G*:�\(4TOB׈&J�pR;��4Y���觟F���u���ݝK�ꆅ�"0�oH�5G��tR'w��5�8a�j�#'8��f<Ӊ=�#H��gG_�=sR��yp�0%e��Yx�C�����"h�Lx��;����>�jZ�j�&��Y�o� \7��S�M�j=_P�ňəFg��
��*
=�=h�����i-�4�N��埖_�ldLt��-Ǫs��Ň��f�-�e)@���Ϸ�\Q�S�]�Q����8��� P2P�T�T,�JYG��WEp�҅��uBҌ>V��aÙ���߽s�����qe��Ti����x�(0�7k饥*9�Bg��z+H4V>w|V
���ߞ�VaG$�������1�*��r���i,l��Ov����f���=�g�m��!&p"�$���3�4�L{x�$X/��ݚ���f��\�;�p��<�r���+����&\�!:w��Ҍ��^­9�;=�O��z�A�ˮ��a𲶶kNI��h�d^���;�L��i"��]=�A�%�/��h2���ڧ�QR��Ù�3e��o����p��j����d����8�e���Ny�8����%'$�ad�n�6Eⷋ�P׳�����b�̽7H]�es8���ɸɘ8���N�#�^z�����=#$6c�ENDS��ݛ:�W��^���B�>�^+��P�Z4=Y��&�:�mT+J\�_>yi|�};�ҡqF�)�o���99�KId���w�4�Th���;��$*"$��Q�Y�;5�Y�}̛�@��^�iC�WE-(��}M��H�3v����\t��gss�rm+��x�mW/;;��{@牻x9�󍓜k�[ݼ�w}�LzT��(�d9}4���/����Ok�z��]> K;����gd��tJv4��yƗ=���:���ۄޤ��I�{UaBV};�RӒY6�_�q�z���
�@1!�{}���`�NN�iG2V��u��}Ϋ�.�}�ߌ�C���ߢ΂���Ul�i��9�c}����w�k�Vd�l��p��}4-_l�S��+�,��#{ss��P�d"WPɔt��lk�;2�va���������Q/u��]�SS���vl uhR�����6(����|��Vb��/cv}"���G(�1g��_�����\�R|��8�s ��W�/G��u�`{9pL�6W/`@��� ���q��y� 4~{�S?
�һ���Wl�
�=If��m|��/^�K
䚪D,ߺ��V|P�7����	�wU,(J�L�h����Lö���Ļ(q�;�n�͏�r�n^��C���U����I�bϬ,�T�Q��h�=�M%"�#����J0K''f��K%�f���:��Q����!2��"��h�x��{t�����#ƞ����%g�{f��a�/�=%���9/��Ã���w!�eA1KK0KݷO^,�e�Vɝ�F�,ޫ��Y��=�\j�?����R��#����@3�Xܙ�d'Cz�x��O��蓮H�H�niM�s$��ml����m��[�?2(�d���.<|���u�{ts&w�����I{�ް����ݚ�������.aUC�^���]��������5�{c�9����Mj����E�S;�n,���dq}� w@���ٷ{��$s.UT)b��V5���㣝��g���u��sIaN�^�#�;O�#�lt�b��8q���^��m�"�z�'n�����m��$�]���ۣ��0n��9t9�`�Ur��qbw�\j�� z��
x��4����u�����]u�^67E��^G�F#gnS%m���Z�=ng���X�i�3�]r�6&�ٴZJJ*��7��e�ӟw��g����z��S�J�N�,�se^�[낧�5��3�D�%ƞ

�l��5d����ə)i(V7�lqN�C����ͱ�z��-�<8�[We���T�RQJm��x5m�3ة�p1�:���m˿��_b��
9-�V�T�1'<Q�w\R��=�ex�xT>Vi_���ZY��q\+0������LL8�9
a�f��,oFު�I/�� �]�5ċO�����RxR>�4��$�Z�M��i>��_��q�2�9h���~�}
�K
6�+E�*��sw���c�<{�6�K�Ӫr�v4�tU�D�a�L��P찎;���Q�w\R�����׋<s&�_�o�lc�ϵ
�8P-��{kӝĸ���s&�v '��ZX��������ߣ4��?$�W��Ȫ7h٨T元)�A,�g)�^6��C�Ļ�4�^�6�m�e����>��w�}mV��l����O{���?�v`�dml�3"@�Ta&t�b^>�h�1�H�JڕV�(L�U�g�=�4���}�W}�UX�u�Q��$X�as��� ���h�8#f+Xu�sa[�ͼZfҳ��'#0��N�l��y7#����d��3��j��Ȭ������h/ ��t6;��;��>��q���o7Ď��8x�ݡ��U�\[�)�Ez�	ؽ���3�'���H�Q��n)af	ݲ�rf>C|`��!��d�f%W�ZI�5�Z(<P��6�a$��lL#��ic);k�+F�ad���a>ĺ"aEQII�d�M#��euo��xKg������m�*�,9�
�ͺ�Ϗ��'_�B�mX% f������Z����4C	]�5��O�u�YIA⏽�qK0K�]��8��@�T�O�x�ն85ys���5��H��J^^nv[��(��A�B��j� <��Ǭs���Z%��[5���S�M̗�����_0��x���m��~�Ud��W#�z����o�M̒t�(v�M���5V�x_�7^��we��Gu�L9&R��hg���c߾�f��|5���L��!��܈��?4D�Wؾ�ut�W,F�LSG�\\o[ވ�~�Is��~y��SEw|]��$��fr.FK"ϭÃ�7Y�uwT��r�\�4W9��K�}sޚl��6ܞ�ĈWP�9w�L��+�.��N���D�2������n����Ͻ<�xh�{�I�ķ��U&��Ƨkײ��<7<��"�0/��i�\8��%��Ǩ�<.-����y�-����X��ƔI�g)=92k��*�8FUMdSNM ���lڹ%�ۭ��[�c ���EI�׳f�\Hbaݮ�Ӭ]o�q�W�$r��X�~]�	5l�f~����MA��ʧx�D����馪O��gpGi���%��4��=z1�Qzd�]w3T�����o2O]e]Fg��H�7=��馄��%���L��ZU�\T9�m8v�&�!f����ݻʱ#4T<w�2�P�����*���C(�.��M�
�(ϵ��ׯ�ˍ�e�T�UA��s�ct�usř�]�{3�Y��7�v��>�Cu�fM��c��5�u��Qҡ�vy�P��_�H��iK=�sPF
G��:�^����;piK��2n�Mb��|t��΄j��V�n$ct��,���}ʫz�*0Q�yVvJ��<�Ԏt�ͼ�"b+vQ[@�Ю'VE�Wx3"�f�#3��RxcT�ʓ�ȣ׺����3�^ȿe�9rv�a��;:�4C��Mj�P=�^����;u�8��g�˹�~�]������\2M{�:�����$mY�*]�ߪ�=~����V�Mkl�&��6�x�cqs�Ӆ�	����n�	��+�aF����TE�\D�z��b��#']�)ċ���n���U����EVظ.���ם}ӒG��vU�����/| �uqr�g���)�	�X�{��Z��Ə#�l=�=���Y�}RWOĳx��n�ւ�P��3|�9���oL�����a�܁��Ә�X\SjAp�����8��<ub��~�C)cdk9IO�N���e�.�gO�2��{�� [�
�����I��p��x4��4���{N�{���m^�N����0X�&3�hZ|�ng 9�ۮ���{��,�z�/���l2���@n&|�-+s^��&&ݐM�'�z8�����]��A�5��k���)3��I�Ʊa����9�I��|1O�k�y�OU��װ�m�0�lg���Fh�ۑTܧ1�� ��o��ܚ���`�ð�Y�O7G�T�Ί����oo��w{�{�p�X��u�|Ƿ��6�g5�<<�Q� ��P��*���.��vd��1/aF4X������w�B�s7�аreПWC5����G7��/���NN�%�h�i�� �e�Z|�w�Ӷ���<�U�OK�mε>�s�i�|����ޙ��^>��r����,a9�P�g����"D��0 J�2!�{;@���m�����F��L����T����e�'r��1��{Y�v묃�.��&�|vg����$'�κ<8��<��N���lF���^���X��|UP��l��uWHeҨ����w�sL����.(	:h��Zb%�0�����?a;,�����c���X%���[4�Px�l;��6xm$�溽�����7%���ο�C�3����d:�_{�II���o��W�:��{k��֯��Z����ݒ�����K���3���k�U�5(�j"ʇ&�`w�i����I����`+%"Ϛ]��W=h��G�w�m,�F��׮fP���%FewMib���eD'v��0�(q���sğ{v��L� �7��� l����K	=�W��[�������f!D:�����K��ⴱ���͚�NfBX�����s	�9�u��'�rElnN��� �=�$��!x��8������^�Px�6oh0Yu�>��Jӌ���s����Q	�l}����FI��Gq��*2|2����P���J#�|[��t������=�E���*4cR���M�13X�bW��sL�wx�����;{7b�s)Z�.Ӫ�2�����%�:#^8��F�&���H��;�� �w�Mf{OY���(6봀��\��w�bNx��"�H����	gu���g�c�ު�,$�JsP���B:	�}��-�s=5����D^5��9C�����ml�@瘗���U�1F(�U
��y����%��>�sJ҄�Y9��ɑ��������4�����ݰ��m�N�\�%��[̓���,�xOy��-,|�ح(}��m9$�!���[rѯ)]VH��3δ���g�q�o�z�~fP�[�fl�M/�<%�맬>{z��9����l4DR�q��i)tTf��³
w:��,^�ߞ��.d�� j2�zk����GJyqD/$���RPx��٥,$�����ճʗ`������}�׬(�ߺ�=��|��GJ�����X*e\Ўn�{ObE��]78��̣�9W�ڼ�j��y_s���	b�VIK��#�1��[�IPIA7_�źK	֙�mLa��Q�v7;�B��{Z�Һ�rk>�\`ޱ��t}۱��\]�v��>r�F6��϶v�ѻ^ު4�y�t���
R܇;TTR3���uځlv��#�tz��\v��G��\y�VϏ5���a�T"�ƪ�Kn8^;9�ݻmk��xWz��͗����ĘUÌ��ewIcc�8�����v�;�;��+ȅ#���_/��u^�Mb*�i�b~�U���&l�����k�X�v�qo�W{9W��Q�鳃��{/T厳v���T�9�Œ���i݃t7�W4�JC��￣�-���݊t��%�i��ŋb�UaR{ջ5�����~3!�!(wus����,$%���)��gH���&����'ZQ��q\+0��s�, ��>�Ҵ��n��B_�oD�2�^ħQ/\+����,|�ץ�����!![��5Ę+2����.?�s���[�@���KI�k�i/�BH:뺛�4�tWiX@���n�abÙ��! ������I�N. �AT+Qa@�ևƖ�߲g�m��I;/����jĴ�w��Vx��3q.:��k�/E�$�V9ar�J�z>�ɟls �mrlcY\�Pu�{'nx�u���s�m7n�
�)���x����� l>2��i'<X��ҹ$,(N.������<�ƾe���+P�%12��l��L�}�V�
�]`G�x�.dUZN#Z/ݙJn��ֻhtdd���t��#��nef�@�B��@�l���:�
>e�ě#�`�$�c ��[���t�؎"N��lՀ����U��'�0@�C�7��r^ �A���
4�lV�^ JM�ߞ��͉�ŧ���;�����`�LJ>1��=qu����z��L�� F:�}�r������qZ/��9�7�mr
6KDh`b\q�yiB�h�Q}�e	AݑX@�zs"Rs�S!J-�35�q'�Gq�֞$@'�h��U����ob�e�rd�@=��Z(0�����s
�޽aRyio��="q�9Zh@6�9U�&���9�/`.0��0��ƭ mE,Q}��i)��ըx�t�q<D�V�-,��)9�Od�f�I0K۷O\�3;8ƿ��#{�4��8���rJ8�l$�\�_=�̼ݤ��3��2�q*4�}S�W��=��Z@���ݹ������aK���K؝^j�)(����ևƵ�gpδ="��R�L��L/�������$�q!�]�S���*{�]v�EՌ�]I���p��3/~����.+�W���3�-5��lEC�K�&7ji�]���1{�#�\(�<;��S�'}	�$ �H�pT%{�<�� z�Y=�Z�&���\�Kҡ't��ԙqF��Gn�/F^=��{��6x�ܳXE�4y;��|x�8}Gb1����1��I805��z�H��8��)(<I���)af��N2�8��=�+'����$q��<��`�{+n+Eg��dà��&�z��,S��+J�۷��u�<~��K��ږ�T���r�"휡6��G��=��|r�mc�B<ٞ'��K��\�#U�h��(bQ����<\c���n�����ҹ$- KK6;<g����I�ԷڄP+��믅����׹�:��`J���=q"Ҏ�7礠�&f��,9�-vjwd�ko�T#�u�X�K�c�_=�}�8���;qZ+�BB Kw�Iq&�[���4�o\�"��X����,Y̘u�%���t�NaC�g*XA�].xW:e��EJ������9�m��wh��4E��V9�F��(z����!�+��R�}���;�]��E��+:�w�Ȣ�	��Dd�7(YU��N&�s����8g���n���XZgJF��-0$5o]��G��=���X��nfފzPz��p;�X� ��G��K����a�r%L��!*�Px���i�s
9���05�}Q\@����=a"�/^�9�_��Ӟ�:�mn�8�R�m@�lpU����<u����F���/U�zt9��������~v��m����ɋ��^���^����~�X%��;[5�°aΨ�H��?�U��{�)���u�9@y׏J�en�i̐͂ eB�����I9���T���kjkNd��$`�3W;���@� �W����wJ�A����iG&�t$-��5�$JN�ߞ�	{�"4@DL��Y�I)(=ɚc�8��gw_���xK��b�A�Y���kXs$(BB)����^h{x��u�%�[)�q���^�ߞ��)��;@=��Eqb����� �4c��Ȓ� ���g+"�M���QQїUϬA@m���[+w#nyvPVfs����t EK�ؘ٭�؆�e�������[6��Y�|�L@���h���/e��o.���`�]����ݧY�7cMM�cG8��oO:���ܣ8��R[y%�̈́݊��
K�.����v��4mi���I��i�k&�G�q�ٴ������k��q��6��F�\KƱ�`wO�1v�s�]vy�+���X�vx��\�՟\���u�y�m�Wq���+���x��Ho幻]��@E2���X&t��V	�����'%�D6���j�G��"K@�Ow���{p��Ɂ���뾐pk����_���Z�L�S��7<�{��^hz\Z���u�+�Ÿ���=]x88����ܜ�h��>k�	ac�ֽh��C����L��� .$�����k��s��O1q�eD�K�,(�Ҿznd��  d�aGn�E-(��mN�a�g�/f��L'�q�6�:�\��DC�K913\)<Q1�Ԗa��=ig3!'a����oz+��eul�NxV}�xB-�Ș"%�a&s3:tP3uOq\A���]ҫ���k^�Px�en��#����4T/SI���?'��Q1Z@���z��
�x���������
;w�)aF��z�g�g$џ�w������Sv�� ��mlq�^u�=�;�ҽ���ܮt��A�7R?;����ێ~���⢶Z,��׏��u���Ü:��,S��+�0���ľ=�}ŋO�8����)���	�W�>��b{:�&f��F����*�����&tE�Q}���t`���dYBfB���o2T�H�MN�Y��'km�ŠuQd���N��*V.�,uP�c2�;�f
3D˗��v�l���6жWxr�.�Jy�������}���"���e��v�wa��x|�f]W�����^�}����#wJ�2�ِM�~U����Ael�AC5�>����+Č���ج(�c�/��t���%&n�tR���P�ԨtJ�;�IXY㙭�	|N��W�ZH��ʴRx�jwi-Ù���������_>�[�G%�pn��_�afF^�%'�9���{�K�>�xVyFo�X%��̗.�~�pxx��=5����ًv|�&ϥ��x��=r�ͺ0�vzn�=����8�z��V�߳���jw����ֽaVnVlW2c��K�+{貒�
7�8<<l� Q[
\\x���s��֔ZK��_����h��vUj�,ڝ�Kd�o6�>���~rd~��2 �+ y׍+=��5�6+5RO�.j�[u=qz�C��!;�Z�^d�Q3���*��s���YW��]n�$tGp�}����8�9UJ���<�oE1��[�&�.���f�ʢ�\�����Y>��L���Eݦ8V/{�ý��Pl4Eg�w�ZA�)cWf�>�*Ï��mn��L��N}�����Y;:��
����ei\Dn��,�K�֒�U��Kd�WEp��oSiF,�ߦ����2�v���K=�i�xNK��H�fb����Z����L8�}Eaf
����KFn��xTx���w�P�g^�׶t*��#f� <u�A4��:o�"B �jGSҟ~kM�̒���Q�LLD��X��ܫJ��e�V�,,��ҹ��  ����zޖ�`��{5�婻k*�m׶�kxs��9�;�$	i�#���Y��ަ��,S�[�31#0%��Zt'w!K�N
"&b��ifA��RRx�ٕ�KJ92Z쁐�����,�Y1�ʰK��
��	Q1$��h��33�|M�RZ9����XX��{ob��a��{"������Y�F�ͫ��}n�t����ҵ����J��O�p.=�(𚝴���;U�+vj�w��:�
�=�YE"i�J]:��YH��p��FfF�'<0٣��.*�t���;{��{��Jѹ�g� U�_"�>���6����mYI9��K�$�V+T(L\u�ӧfu׶���Q~B@̲��*�KJz�+E�+6�J��5������2�B7j���6��G��:�.ݣ;"V۲��gxy��7���|x<4�d���e����C�s���5����b�s���W&X�7:
 K;����d�#�Ahx R�;�3*�K3gnkNLĉ�'0����-҅>�ⴡ+>���ĭe�KD�Nyϳ���A��#���|9���I0Kf7J�d��%b�9�N���KO�w��gZ�����':��,UQLm$�d�� H@���]⸡)7���>,ߢ���34� d�*7��1y�m.��߾�+qR� <���v�V	a<�a 2��zk�N�W;a&
};���+>d��������ª�|���~h������0+Ղ-�]�OW�xH�g),�P[�-�lx�n_l�����:�"���������\�"��^�p��3u��zU�3��F��O�{�%��ӹ����^M����`+��_J�=��^�}����O���7˽��u�c��P��M�:��;�!�1��tTq���.����z�+���$����$ҳ��y�ݘ��S���d�t��I�Jf��܀���5�Ǫ�J��8:�\�1կA讕[�`9Ј�l�mS�xz�ڋ�x�;q٪�V��u�s]CU�y6�6t�9�Mh;�Jwch0j���C`��q�#4^Ӝ���ǃX���]�b�ޮ��͞�QQ����m�r�XVWQs��"��`1��-r�e��+����H���4���^i^�|.FLB�h1!	�}4e
0T�1W2���4SfC�&�#���{��w�+����N���zt�݌ ��"���n�������u��t�r����NK�b�{�R ��ɷX���ږ��V4hȝ���^�����F|�rN���ٷ
B�u��H�>]Zol�b6�\�nb2�8���1��l�j��G^,�':it�v���X1�1&Ч7.�
s��O�!hCj��ιU����2��������Kʰ���,"����8e��"�;L��ݱ��UR����q�RF��:b&��Cm���D�y���e�Sр���b��킠Rsn�˧���Ie�\��o�&z�;J�w��h't�;�o��J˳��L�;�h򻴾��P��/]�W.��s��u��Z��WA2��ͺ�>��)��9�v��ax}�Edf�	:�z�ۣ���o5[�9Ξ���GB��\��;c����'=��YN�IC�q݁׷����odcM��͋�xl������hVL#����<���K����"���ו�Z�5�\q��ln�oF�y4�<�uWo9��90�&c���u�`q�٬��m���A뗱��ggm���[�>�VT��.k��^%q�\b��׌r3�wS�n�[���uʹ=�:�����T�ϵ�H�g+���v{r!�F�:͜'1`sv�fꌇm�;��:��]�X�^�u�͕�5��	T�m����vq�T��y����,��Ʈ#
�bg���IcG4��7U�����Ʒ-uQ�UV��;D���y�k�8\gaт:wcOJ=q����x��ND��s��nr�Et͢s=��[����y��gV��u�aH�{N�&(!��3�`����"m������l��<kC�}��3K�黍F���ǭv��Jq�ͽ�nz�gSVV�v
�P� H�65S+*ݴv�vg�&p�4`y���97WIr�;�i6����(��y�Įɛm-���95֪��: ;�v�5�o5���,�����Ǟ�s���ss����.��{V�r��X9��z��v�rmI�ٺ��^ޝq� �j��2u��y����۴cJr۞�yGeۙ�y뱞�`qax�{]�������b����q�O�`#��^���f��ε��7nn��S�:)�c4+�ݘ�rj��m��r�[{]�eͷ�v�ik=)��nxT7��i��uZ��ю�:p�Y�$N��fѸ�x��p)�f{q(v1�u=ڑvK�s�ۋtp+��{���}vq�%t{f�d�`b��`��H&h��cb5*-�A���3�ےy���8b��c����]v����x�h��e�M���ц�q�T�1�n5��޷/S��\�b��L�n��z�X��lB��o ��s����.�8�cv�vySR��S�CZy����;���[�����j��!���'X
YU"!8*��z�*�Tƛ�Q�p2i�Xtp�0x%]�SW}��iIP�5^��R&Bji�S=�����}���g�͈��Z��c8�ޖb�3on�	��<�N�q;�C/�G���4�\�����ݾΊ��0�t�G��힪j��^����5�ҍ?A=���S^�*�������ry=$#$��g�h;r���q���T؂�{��B�u;�ѧ�>�nS谹�_5�9�+ُ�<wū�{�:��cڸ6�=��O1��Wzn��k���q�T�.I� �x׌�S^n��uːl�u�`�E��^\b9�mͪ3�s�[9��ni�,�����r��Я��K�"W�OZ�!��OXKۺ`WNPI�AjL&��p8�x��x���>��M�+�����<�`@���Sʢ*�r�Շ.ҍ�g#��y�Jk�����������
{���t�D��,�@��Ē��ې�eQޏ��ׁ�0�m��!�쓾Dvzr�����<���uvʷ��@�������l�h�y�����}�2��l��YY	����z�����������en����P�Q���\%pY�[f.��Y��uʱR�5��vC��)�pu��N�z��9UL���q��о��}��GX�r�u�77��&jA��(�xq?:�[0/87P�G�Zq!"<�n� S&ú�z��k����+�;��h��i��Gvi���\�ﺒ�h��h$���c$��2x�k8�-cv�'����(�Ǟ:�ѫv^T�ö�vyU��X�����;M�.P�Ȋ�n��׶yo�&�;s�a�i&۷�vf�������Z싱˳�.s�ׯd��݌�K;���%�Uٗ���d�Sh*]a���3��=��rJ��90pq�;��;�n�{ e�v��[�Ⱥv� /K�C�:��u�\��Q�lj:�*���˗�r�[���.�G�q�@�8�g�w�z{���S�#,�x�����>�s���1x%ǳ&M[)�x��r�2�p4�1\[.NŤ�n{a�n���]�a�7W\�n�Z9��i�Y3S�8�T�Mȉ��b����))<X���- �-��U̘e ���|du���tei
 D���&&e�Eg�3/n�y�;xJFe��?dW��{o^��aC���1/$�҉����j�
��F�����\Q�Q�����ުѹ2�����:�f��,S�Pj�N�Y,�={Z�Q=&�k���ŋK'�\���,|��KH0�a��HuF� �Y�ܪQ�;�(�&"eV	a#�ֽ`��G&d38�����M,]Y�W��r�b��ag$�w�s�)=~�|��l8��x�t[=��=���s��E�9�4[r*�cZN3�!)Z�LL2�,����P�E�5��l�sw�z�drC KK;��+>�j��e�%��5�>?�n���o;��@�l!I��3����1��D �zQ�����N$S��M2�K3�4i�����8A��,����A��0�	⯫=;��y"���P���у�*٥�n�����m��>=�r����H��:`+A�`4���C`M�q)#�^�X��k+U%�=��aɘZ0 J������\gq1%q
ɏw:����v޴Sɨhd�@��9��]7ib�ݷ�%ffmH�xA/V,�f�	����IA����4���9����9��	/����<-����D4LLV�N>m�a&�00$�|�
�ٷ�XX��}9�%'�<���=�)![Em-uB��Y�9��#�$ֹsn�79�e׷GK��w�~v�߁O����ʥ�	GF� �=�{*�K
ٶ�ɚm�I�}t�Y��p^i�쑲;Tn��u�����g_��0L|�Ok�I�,��ץ�%�nm�i5�>5�ں�_����!����h��v�lV�NdV�a'�����_a�A��ϧ�wIj��Rb�6��U�镑��/�
0�N��d��=�b�I��"5��;��I�Gn��Au��᤟\$2^ʰڷ�x��13+��8n�~Q�͋c�4LJI�+��uz��{_�"�ng�H��`��J��I�1��R�P~A>F�]8�i��޾�f�f��$uypP���bf(	=̙�H�>7��R�O	t�i^ �����,9$���;���Q�5=ľDp����k��<k���ͱ��M�
}��iB��c��I9��ݭ|]u���ᨽ��TT) �oj��{n�0d�,�{!�t�	TۍD�#L-�>����j�Er�p&q����{��3�.1��lV�O�+]s$%�i�
���4��y���KMY`ο����n��s&�L�af�u�-$�.��z�'�g�oeVɐ� h���b�N�R�	�	�&+EG�6���I0�<�j� ��N�L��v�\P����X�{>��]��vIA��\]a��'fN2�������	a&�W*�Ҿ����]W}��ȅ ��}E��:b��sy�U��:a�K�D�M�G�D^D��.�fc�l�Q]t'��"���Q�Mh�pV��L��2�Pj�^����Aذ}�:�[�}̜��ڤ/pGL����:�����\��ڊ���qgwg`�����I �	�E�Ӄ|I��N,�C��D��"bf�X��z�b��a�&d�8��餠����zZA�[9:�I<+9$�N��?�{�ev��#N�u�t�AH���:�9z�/%�(0�B�)"�k�鵤f}/�����Yh��X�}�q����s�ci&,�����L�%��Q���\X��{��b�?�q�(;m*ć���9����I�D���]�=�+{~+��vkb�]Bd�$c�X�{P���*f�r
L2k�}���<�Ɛ�o9ۚYɁ0� `m0��⒓��R�L3�Q*1
x����2CX�02���s��KJ=�����Y[M��s$37�ⴁ*#��l8�@r���U��
'2�%'�9$�jFm�M.$�K�����±�w�K��9n���RyoZ�KY�w9
��;���\�ܲ&���G�E8ЄGc��6cU��T�*�Q}�*��\��g�۸�ۯj��Q@������g��.�z�g��6�]q�p�v�p/r݅��#!��$��۵�kV�����Y�����x�w7HN�/L�<��9��s��cq�b�㴻6:�<O
��y�nۂ�cK������`�w[^�M���ni�"e�6�7Vw��v�3�OWf�ք�f�6g<��N�%.-ԡX�4�@��d4I"����
�r��
K�����修��@�G�5w���[؇[ޙ�>�Z$�Hn��4t�@ :��k�|�]��O�{�d
��r���<)��K\=�h�6.0g�y��8YRv�v���pb��TU�Fʉo�����V�UB��0�h}3|�ٮ1��h�ެ�ƕ�no�\�� 	q�i�;u�II����r=vUd �b믍.�;3��OB@��*0_���%���z�Y⌭��ә1�M<)��:
"�N2V%Gz�����[oIO̗&hM"���T�$�K��,k=>C�C��興���gP 0j7g~��I���S�a&
};����$��&_����?����v���Ԃ�$�H���c�ii&�!$�%ճʸ�gF���ۊ�I�L���P� �_-�_��qN;HWS����A�8V�l�;�G����k�Ԣ�O�B�
��v�7ib�Ҽ@���+
O�lU�0�_�Ƴ�u�-(�,��#�DP%)3o綾{�s�s��g����^��^�2�E��.l���j2�{Vx�]��c=�t�~��m#�<K�u�j#'6e��oH�b�R�6�q�o�����q��|1�J�<�W����
�ɛ໨���y�.|�^��!ė(�^��=W*�35f����R���kb�PaD��l6a�Ӻ�fa�� d	|b�ޙu3w	�&"������u�%'�w5R�I	h�2����0VdWG�XX�9�k�M�i�)s�W�kZ��i6��w}}MÚP��m�ĉQ�����aɓ֗C㾋����יTJ�^�e�i&	F��׈</�2u��BK���U�i��=q^�(�ݛ0�v���X�]m��DR(ڈoEv����be�yz�ܓ�Gm$���l�G����c�Q��R�8���s�����9�IA���n��d4��A]1�W`�o �����<ˠ�����ͭ�ә0�I���WSqf�.��+	�7/Ua̐����|(>-P�R8�U�!5�WǏ~�x�׏�.��fN��hdN}ّ���׫�J��6A(�������<÷Lk+�K#6\�&ފ7�f�ʔ���
�gz|H�DT듈�opȴ~N��jɜ>�躤�͹|�k¼�{�����׈X���z��-����Ī���Z(9����3!�m*�REKpO�3�u\�y�|<9������+�,$�ڸ�(��D�,�\Ǯ:��j%��z[j���Ĥ��y�J�[��9�
D�|uos��	��w�Ԏ�
"%�
<*7$�z�,+�3�i��ޞ��A��M�|-��U�	Q�%ۮ�Cw�06�mǮ�KvYm�[��>/	��t�t���.{M5�ߝ�~�ϯ��ODD��E�;��s��������6���2R��%�����	i$v��qD���"���(�ʝ9�����0WSܫJ��o}��
22�i.fa'C$ ��|>'9��x�T�ʈNL��.(�.�ۊ�O
��+^�nfBI��|>�tV�(���m ��Nw*���4���Y�=ykOQ�4ց5���*�E�պ*I�{r�iiC8��*!Κe��{A��VK�<�@D"ť�6�;(k��(��H��89`4�E�B���x^-��S�#z�����p��U��YPs.�P�Rs3����zo�̠.�O�L� MطZ�W�b ���) ���m�p
��/!��*T�"����	��>���]�"��	\J&�%BS1X%���W������U���I�N�XP��{7�,XQ�6����sp����t�;]��'�m�Ŷvx0�&;&�q�j�����њ*�%RD��%&>����L�ٸ�(�����rL3%�ZP���Z(0�`�/��&f	O/$D�iF-��+9�vT2��+7��U��J'0�zJO{r�iq�i�k�~q��k��H�n!z���,�|?����,$�ڸ�s3��V�u�i&����^,JON�<�GE0�ο�疗jM4�I���]����
w9�i&	l��֒x䐬d�|vߟ��KJ=�����C��`��G�oi��
9��n�/�i"TvV�XP�Y>Ŷ���,�r,�����Hﾜ�iդU|2*���-R�~�Y��Ո�Y90̋�����2}N��B���`�'��c�L��y�~G�Ѻ��b֨.w�k�{8ݽ��χQz��n1����z�+v!��Er/���[t�\�w4�l�=�;���'����':M\m˭��ܵٸgq��1�oY����r
�<-�=�vAe;=��bn۷5�/s���cc�7�-�Hݰ剗n�񃉃�^���^��N�8����v�<-�f�mdF]&�Il6�H���G�5�lf!42b"��*L��^=��_�・o���.�FO�ߗM�{�o�U�]�<���8��Q�6n�mC���F��(6� �x/Wa*%��%����G���;r�,���p��iu���5�$Q�p�ŷ��K�碴��Y�}���=�V��<@G�JoZ�_�c;۞��_�s��$��a�bUaBV}��=iɐ�/����ފJL$}�qKI0J76�Ӓit��T`�oƉ�P�0�Dʑ��	ic�V�h��G�oi���0��fKO��Ur�$J��U��
5�\�!�RD@��IIQ�ft��^7z����]1�W�<+s~z�,9�@�d�!wu}s�c���a:���QHZ�S0ɮ1��S�Uℯ�3��ٽ�,ZP���II��f�������_<�,� n4{Nl�.u��]�u�c��;w�T�f�¼�� �������	XE%q��f<��~�����kb�Px��u��&B_�񧅽u�֐%Don�<8�C�B����c\x��y�h�v���Nz|A��jj����f5Ii�\�A��C\��B�{*�N�x8��"V͕}zi��=��$�! �i��uD(1�]�s���O�=���U��;�!TT{pZ�f�P�$�\I'Hz���X��b�&�Uy�漈w�v�:�3+�z��I̖	��+4���qKĘ%�ݢ�Y�|<�5�fa�HO��F����1nRg�3ܾ�k�|
};��Q��$�$�7{�������{x�w]��iu@R��Px����L�&e����`�ȧ�z�,,}�׭9�	��7��n,���ۇ��$�4�!���Q��Ұ�a|��}vM/�y�(0��:▔`��mEx�³��?���E�n�x����D�S�h掮��[��=�p�CK�
��ۺ]������$��)D!D��h��?w[֊ONdm�i&
};���ft� `L��q/�޾��u�8q�T8�ݎ	؈��ݚ[�3�с���Ļ{�z���}���F핢�]�/� z�'�(��br��8��h�ά�/��|)�0</������᜔"Ǝz｜}�=���"8���U
`�z�T�%�R6�{����ٙz7`��OH��pf� rzo���������q�iޡ��2f&���\]�h4ČK{8=�(8��6�W�q�{o�Iяn���X�x$f��Q9�Q2��U��V`��݈1[�hyIڗ@8wv��P�{bΡ�6<�x$����X6�ո����M1б��Zn��}�0z{Ey߶�|yJ.[���\(�]g�Ng�t=�����d��h�����t�5�`�7�3��`I�l��A�&�LU��.=T�ʮ���O]f���f�C�6yS��8����B�U>+�_�{�ɋs�N~��$�SU��ᷳW�!U@�v����eOw��?wj��YW����ڦ"0ų�n>��s"���lӺE��ë�ćs��#�#�sΩ9�-�P�]���c��j2y�]v���B�����%в�����|������Y�c�����4s�W�������'g�]��ǆ'�.�̛S�w�3X5�h3�ν�;k��P�ݚ*�D���8�yk0��o9�/��N�^�;}��L�M�<���/%�f<��	!t_(����K?�W7���p��O�2���{�1s]�v�z�G�<�Ҏ�S%�0�����´5�(���ǔv�LZ�<��'!9A��L��?췾=�2���ߥ#&���C}�� ^�yP���c��x7�{t{|�m��#��%����3�OP������J"Ⲉ��ݶ:+���'2����*HFg�h����b*0E���w���=d�@��5����H�1���gE�dj؍�u[b�T�w�4�&�%��W��Y�t��|6��w�0	ܣ�m��'���:��o�G���cW��$L8�n���7��7��5�0b���h�
hl`J��̷�7���������\�:$�M��LT���\���3tIoyq>��=w��AW�s|�'�����T�20�wm,ݰ]Ƽ���fK���*�!�����;��O�l�����6f������(�3�כ���?�oa�/C6�qQ	�6�����>��n�nh�qvu�G���e���Yk����0kÄ�5[�I��{Q�Ux�u�J���c]�d犕������48R	v���C���!�����T��K���>��������p���艺.��mS�s��/���<p�zo��u.����@	:��7{���^����N��e���q��I^K�{a���Z1,�N������?r���s�2����ɽ��U�A��]�}��]8�gZL�]�7[�2{��<����
b��n����^�Pw���׵{ҝ�7;��*b���@�����������L���'�a"k���t��x}�g��t���[�]Ѭ�Z�Nj[�Ȼ��H�c&�Q�������m-��Ke,ft��Y����X���?_Sfpˀ�1���]y�?Ku��g�/F����޸�\��^�`����u8�������c�^��4)����N�tM�B�0�e��KD��jkEII�f���-$�#�uje<���L���׈<rLX����WvM|%��ݶ�����n�I�$�fKmg=��q�K�ż��C�ښ�E�����
3/ni*<Y�0� ���iiG�]�����Q��X%��.�\�����t�G\�����n:�p-�6���13���V�
*�J���ޔM\�-_��wfF��+�g��M��X���V�%F�f�s$3%�O���I�,���5U-Ӓ��>4�{���%�f�`�F�7��%�[5�A⇜ݤ��e�2q02&����\<���)@�/2������,XY��\RS̒�I��afFwM-(�ON�k�m|��}�8F��Kk��I�is�$�̾2w�z�Y��M��P�g5V4�Ϲ�uw'�	�I�"�s�׈�-��Ys�{������������'L�Ϫ15��	S�w��ЫR!�wܼ�u+�����܇��V�ZFt�g��mRo�8�qa��n��g�+@����{Ә�KEM���S�w��!�]d��*e�~	��d
����+�J�O�4�y!9�%�(<I���KH0nd�$�%���XA��#���L����A���.��o��I<45bbP�	�Y�	misJ�X��+S�U�7u�V��{ߣ����tZ5�2�0��P�I�Or�%g�of��aF���\��Fdgt�ҍ7,�yrZ$��^%�H<+3$ߞ��d2g������PaGWV�h�)��U㵤��������k���$��J�5������(<I���KI9�%��븭 �Q����	a$n��R��(�O35��ܓ;3@�Mn��X����I�[�iÓ0���>/��zJ,�r�VA���&f)aF	n��V�xW̙�/�	�-�=�V%���������iF#�5y9�/��3�ܖ����F`G'�{p����HqG��&����ͱ��3n��i�W���E�����bj,�֧3�+5�>N�9��po^8�=y�#���ݛ��.�l������;���`����[���kt��m�EM�R\6w�fy@�tc\v7jkǶ��agp�RF���p�k�^.'�s�sXrv�ۋ��N��J�X���W��\;tltS�61c��_P��P�9�nx�3=ػV��u�rllqY���9Es֐w�n�g��R���ǑG������al���y�z.����'}��ѕ���Ó���t}g�f>�{��|sh�����t�H@��-�������@\5��<W���}��'��m�����k�^�[Ek/AC�����Ǉ�iD�D#&fEqD
-��l�p��zI�nmlW30�IqD	s�s�:��2��MU�\���q��>F��i��$�
� z��K�4�O��V�%g���+Nd�ɰH�������%n1��m�ī����޸������I����X/꣊�KK;y��X��ͷ��eX��P�J3�'�2M�_M�$J��oMab���V���9�K�xI�~���. �OjyT�V'�$�m����w��g\'�'IH�3c�[}U5
&7z��>�wUiBVre��y��@�Ԡt�m����p+�<������*�G���7]:u(�����Z'�/ѐ��e�J<�k�������C�۱K
0Kgv��&(�9��|mj�z�G�*��p��P�S"��1����]��)�;�C�_(��Z�k̬�{t�1�F���U:��F<�q�B3:�;�'�P�#�̌��P������c�Q ��M�bx�t�D��8�e�ue[�����R���H$#f4��9�S׊k#$�кQ�k]j'6��� ��	�h���)�@��O����+�q�>8��oU��|�����X�\��`�<��
�F��X730�x�%��w5
:�����,Y�N�F̧y�!;��3*�����d�K�7�� ZQջoIA�G�f�aɘIL�-z�ߦy��|�rLn/V�l�Э:�,,|ݸ��(�I�d�4f���Q�
v{b��+=>ݚ҅��$�-���w�=��6��̌k	�.یoX8�Ǡ������`Tnt~y;�;ǯ��v��0�]�D�%v�\RҌ��j�xTz7~��f��-(���Q>R�O&��$K�>?��ug}�|҄�q �8�ǳ{"��aGn�qII�G�f���:q$�K���S�C�;C�<̽q
ͬ�uX%��������?��Z��j"�d���_7/t���g�^�qƺ=� �7�rr�-���og�@��Ck��Un��g�&�4�Z�.���H�ǆ�k�b5޷w'eU�k[�W���ޔ'�i���؂`44L^9qQ=@
�,D�����>���I���}���������gs�:�K6�,��U�$`���ab�L�� XOJ�=%n�tR�LםҰ��&HL����Eh��mw#��O�dL���3�o{��]��a�`̭��W%gw_=a�ۊJs&լ!o@(N�N�}
э�0n�sܙs�tEkמ	�8��-�G���tߝ�w�}�y�u&�m(�v���^/|����̬�uX%����Ɇ�3-�H��k�}5�U�?����:�J��͊Ó!��eb���Z�s;'�)i	{juV̆d���s;O<�e��[��iu��;�h{x�7v���I	7�5�W=�W%dgv�qָ�2���TF��Pp)q(��&vi����T���]1�V�xVfN�ƙ������5X��?m�3Ce���X� \@��Q��w8�NR[ԆQج��o����+�Y]�_�;���}�:\n`v�`7�*�(����ATXE�z|���O����\\9j��swQ�D{�i��P-��{svV�jtΑ�qy�-π@?���f�^3���})P슄)��X����H�L���]����K�w�IA�M��)i	rIJ��c����v&z�	��:qÞ.��$2�(�[K��9���nI��Zց��8�V4+�*�,�|N���V	a񱕪�Rx�cvt_��	��-$�5�ʸ�+<�C�1$��J�w�"J���VV�7&a�'���w*\Q�]1��H<+3'_��%���(%���;�t;�B�D<N�$~��lR/edNjd'MG��L����s��ī��s,j[�Ӥ)t<�R�L��왧��������	a#�f�h��̘o��d]�Ip�-�wh�"%Ɖ���U�	Y{u�
rI�2����J(wr��%�Ƹ��Y���ˣ�zNhQs-<�
6V\�Mm�s�i�s��W1�gq�§� �3��0��_J`�4�]�X̟P�����e��R����	F�F��k\=1E���^�#F�w/h콪�n.���N��8�xծ��΋v�t�끰����x�g��Ӂ�tb�N�EhPDw@�F�@����j�-�ݥ&�����ڵZ/>'��7Q�.ܸ�����n9y���+��ku^�H��)�Zk��y[u���8��A�]&^���-X���c4�����r���]�6��Nh]֕w������@x�#N~;=#���h���0wZN=+<r�y w;�-��x��m���q�����ݢ梖��y�:X�P-�g������0I���N�X�;B��z�n��&���{V�m����]�������eL�W<�Kls}��6*<P����I�
wk^�24ˇ����u�u����~crR��R�=%�63u�o3$�-����ⴃ����+��bsUh��$$�Ky��?��Fh(��LǮ����V�҄�����rd$�	i�^������,(�!B�dC����x�� �̐��H> ��|%���5�I��ݦ��9��X��Ɩ?o�_k�mn�#����5���O�Jrf(`d�[�����,��+<+�{�XQ��g;�g��:�]̛��us�+5��H��@=���z�,��b��|��z�Չ��m�H����Ra���Ԗ�ab�mj�(J�ݽz��2e��K3��zJ�(�Y�P��"�O!&��d��k����=Z����Y5������B��W���~�O�}Kٳr&ۡeo �Hv��*��(��lףы cHH�\X��Tt%������M�5��C�����\�.�$]]x���;�w�g��e�8��p�s��n�o�Đ-鸸�U�m��X|/�}�a^�G�ۊ��FF���rI[���K��s�"b^D�11^ J�ugMa"����⒎d��d��2��z\A�/OO*���x.D��9D�D��8�紵U���Eo³��ݴ�9��}�����$	!&q/�gw���iG���L9J	R�RTx����K
0nd�&q$!7To*�����X%�����Ƿ��K���n�T8*��$��:�܊qkn�����g�
{3V�竰�ڪ7�=�=�_V�Y>@Ymu�*%3^q���vV�%g��f��ac�^�rL�2JL1��ޘ���Kc�c��B��I]EXY�|?��+d�q3igmu�£&;����>�kUi�0�(�/��O;a
���u��?s�������wp���gb��w�i��}�u7bP��\^ԫ�Y�| �p���֞q�Ӝ��kq�;9�=�g�����"Ϡ�H1ϑ!�W@�@Qy�_�=~�<���L}6���e�~[2��AgƬ�x"0H�"���J[�%e�R���.b-s8�@�I͊�%�g{��@fJ�	�D!�DB��D�xR{��ұ@�w���9�j{f�@����U�I��]k[g��k��~�b�jyȅd��K̽-$�-��z�
��;&h��U�ZY�UʴTx�cwi,��s$��G�:'�G��1n{h3Va\����p	lns�A�]���1��zk�%���`��w�SV2eW%fow�XH���Y�%'���U�0͂@���	v��(�Y>9�V��&���8���;�Ϳ%���2Va�w���I�V�iVg�4�9�	$�Z|g|�D?8LBwt)�RRPa'Fg=-$�(��+9&P�,���U�vWYZ*<Y>bq<:י�	��������I�,�_*ℬ����	n^�II�;=��ٗ*�U�Z���gR����6Ep�N��"�WaRDQ���[�qL�ޕKcJ��3�ԙK�@�m!:�`S)�r�%�3�h=��/���<���r ,#j�'P���`���y,B��q@m���1h��.v?��;,���|G��oh�����>P�"�(�D�ʒ��������,'����]�X(0�����s	���i"Ts3v���u���{n-��&=;����&+n��ù�l^n�x���FJ�K�&��iO����J1�U�!�J�ŏ���⒃ě�����wi��!�-(�|<�s։igbд[�u[F�-s�<{u����s�֢�^�4�`���W%g���$XQ���Ľ��IV���u�Q�XK-pyx�T�Q�P��+I</�ͧ���Bq fm(͞���P����J0�fj��Y,2�he&uׯ-i�%��>��t�ic�-��(<I��Җ�a�0��R'd��OZI���n��:9�wQ2��XY����Rx��a���S���9�ur�(JϽ��V,(����? g����y`"�����ܠ�����?�wt��U���Q���~ў�c�s�m�!kq������5���b"�ֹ!t�8�j���ٌ�ʩ�U;jn"���,�|i�;9�[��e=���$ƽ�L�X;�Ÿ��f�̤i�ɝ�Yz�1Wrdw/3}2�iǁn�b�u�O=w6����ɵqT4��J:F�����V+�:�Tь'���O`�ۑ�Nc{� \�����腲lm�͓GGpZ�;1�(]�-��om�3J���u:�n&-+��3ۼ������X��e�>��l'�������ک�}z�|���n�T�����}�qZ���N'G�
�+���:���W\�k{��@D���߯/՗��ζ�մp�$O#(����rd=�oj<#|��_\�����*f퍚�ȗz��dWWb�$�.SYu�0�^DP��
Q1g�9'�9gV5�B�I��vja�Un�QW�����sH�Z��`T���d��A�]�~�͗�2}eu�1�vc��E�*D �f{�QwۖB��9c���߅+ˇ�C�?��v&S�+��{�>�g?@�����s�#� �l��Lpǜl�;S}��Z�������EѬnh�w�V����N�a����]͗�]y�f��c�q�Y�N�N����|�]'ہ�G	�qg�ڿu� ;(7#1��;��̪�_r�v�;�r��t�(j�3_ V:��9+�
��OLF-��J�V��V��p�#L�=qp��i��]�M>ӯ[����<�s�՞ܚ~��&6�rà�r&HKt[J�[&w��'���2XT8�C�6A�듔M%噥��.�|a9�r�h�{�v_"ɐ�.1���gu����\
nN����i�J5��Q�s��f{)3�H���X�<�n�f�#&�1�)3�����Α��Lv�^�nv��m`�M���\c�m�js���v��U�]g�7e���y��2��ݥ:�J�qvC�֐�w�Vn�e�ӌ��z����E�I���CY�+�KM����u8�Җ�ۜ���������9۷<5��{u��{�ֺ�x��.^-�H�0p��q�on�A�a����$��n7[*�uq�u�pΙlͬwR΃���n-�ݻ&�ܘ�]��%����e��єw<�s��f�Fz���%��5�l�{%���[]��=�w�gS'u�v�Gd�"�{�n�. ��N�m�d�nWX:�A��4��a�˽�i��1�n��ڹg�#�g{Z:U��eG���JM���{��Z�+N�u�n��]t-��\�kֹ���pe�WDB�9��<R�&�m��/:/E�����h��h�5zl�N�w;�]J�ZLғ�[*n�]�iz"�-������v�ru�h�^��a{�:ƻ=�U���d�/��gv���]WC�n��"����vݵ�CZu@���:�G]�0�g�mk���f�e��\#�7θNt��^�Y:�c�y�֌�p��<v�,����m���㋉��'<�u��^q��ָ�g�f֊3��'@38�F�����5ֹ�kP���v:�N;�H��r�{fqX���Am��W ����3˗gvv/C���Ʊ4�4���ۋ����mɺ�윋n&6���n��R��ܸ��^Z��l9�㋁=u�;��7\z��u����1�cs؝�=.c�]�/\i�b��s��>w��ݻ7h�|s���&���E����<7&�vr��'���j��V1�D�v��o:c�=���r�g�`�ۣٹ�3Q�u�m<��h���'���GSokp��#�JNUg�Pq[p\�u�����\>
H`��Y�v�.͹gM �w�.��������G-�ś�-������m���t�v��g^P��bD
�G]�����!A;�qs��Z��zae�Yw҂��q����Z:7�~��l8�= �{]~�:�=�u��O3t���C���u�����lA��U2�N4U���a�6HW	T��;��
�;����ӹ�<����Z�����Z:g��m�llM�t�җ�0�EMU�m��6����X�͒�������κ޳�vG��|{1EG'�l�w��G����%��x��	��Wq�=|�^�%;��H���5H=�O��wq��/��*����:n���c�{«����&]CwЄt�t�C<6<�e3J����R曞$u�W�w�Ꞑ�$�U�y5{�It�f�րC�}��o����7̕v��]�9�A)�
��X��ͼ�̧D�Ӗ�
1���M[�㋩�ٱY	8'�����9b��.^�2�wG�0թlX��A�M�:n��a�s�J��|�� r���dfT\4`���3%)�m�C!C�9N^�nE�Ԭ�)AR،�{��Nm�@��9�V E�Ou7,a�)�"������C��W9f��3��>>Og �����;�L��L#W���j�XF��P�!�.��-��u{8M��nǯ�>�u�{���Ӝ�����7.$2�)���[u!۞�扥�vO���?6ze���G,GhHd���V��",j��T���X������s�����`G��cWkF�h����FS��g���vܜ�]�
v��q�v8ܻ��,uH�T��"(J"���陸k�]v���n��G]��t=�l�>p��w8tC�tq��g.ȹ���s��SY���+����n��b�J�wQϒ$昇�cm^s�ڮ��uƳƈ�L��ۼ���ey:�����w��0�U��4(w՜;���x2�����*���+��Hb��
igw<��s	aa2F�8؝�r���ݹ��ǃ���n����������G*n��J,J���y�>	zc4�,�36��2p��-(͞���Q0��8�,�y���Ҍ([�[���H��$�Vn_r�(ZX��|RPx�c3^��Ɇm,L�q�ާ�/�����"�α���+���6��O2Nɖ*����?4o��x���y�A�V�Aơ)3s$�FK�c�褨�΍�zZI�^��+<s2_:X38��+�����c�������&�5���7���Ҍ$��&l����	Q���XP���o]RNx��7�\�����D�u<*�O��_���N���kf9v�d��y��<��'x=�����\����~�ُДv���ǫv�K�ܭUə	�IlH�����$Yף�jfT��YeA(��_=��g�f���R{;>�ٽ�U�>�����.�+a�� I�=W=e��x� l-�&_c����]#};W�b�e��ۺ�I~^�t,F�f�A��\
�(ޠ)b���6n�m�����n��{	�N��Ш��FJ�xY "K17��JM$��ץ��%�Ұ䐚���|ko�my<��r�% �m.��v�V
O>��6�s3/;2m,[���qVl��V�,,�T�tb�%�əS�¤��2N�R2J���z\I�(�z��k6ްKfC2o�����A�=��_1�ҦY-35�_Ѿ�UiBWɒvJͽ��$ZQ�7�IQ���zZI�\�x޹C�C�'O�1!����<N��ܭb�N��qb���u.�nyz?<���<�*�Q�KG�c�_���=h�dn�ׅ'�w6�2a3.$��mOt�%f�[Ds;<(tL��֔,,|��730����Yѷ�K�0K�7J�
�f��XrI	8�@�/��Y��T�O/�"�b^�PaB~���H0�O�uV�W�s��/1��}�v��[��*6X��_o���ݽ��w�z�V�1��s��}�v2Xu5ݶn�y�6qz�N *���	L�-<,�Rv:�Q��o����`|w �N?ZE}�!�9y����s@���!��FT�$:�2$�
�̩͝T)��u��V������5��5ƈf�:�T4f,m�Ԏ�!�䘉�ZI�����d!%��qf�u}�XI인�
��	���#����4�{�T�(r"$�w�z���m�(XW2N��&gK��*J(�N�KJ0J67J������{��QJU,l�P�K!tԜn�j#[��*��kk*�eԪJ�Cp�Z�h>Iu�i2��ϕ�[D�r����.��{=3mW�B}���H0�O�uW&a�f���/Ͼ��L���-�إ�e��Wd��J?�6)o2I�m5�%/��q&��7�Z%�[5��L2T2Ta�5��,AA6�k�>�k|�=sK�=[����$$�H�;�6�<o��%&?������8���
]�Dʭ$�̘L�����g��҇��U�A����6�a]��{���z:�d\���],��a}�u彫z�H+y\��su�8��r:H�3!�4(�@�@m �qYAqY��J����&�G��L��'�F�jׂn�O�Q�\���>Y95��Ӊ�1,����Q�xМ<�Oz�L�}����}^�;V�D멳�φ����D:��W��@`+m���s��e�B�C0$�ӝ����.��U�����E`�rf�돞a�%���b�����h�<��\v�ή�ڰ�y;�;\�v��O�U�q�Q����J�v21W@�
��?)�s
���iVF{uW�0̼2c�Ŧ5��Q�J|�l;�x�*��`���=o34�S$��x���+�Z|?mkׅ�wg���-m�%��澾����#*�Z<�J�oo�XH��s+b��fgL�@�����󷢗xJ��i'��n��I;E:Ք�֗<���KKs���
L(~��m���Z@ܙ�d�7;��u�]x��D�W�Q��!0ī�G��إ��7&BL���V�`��޸�@gt���G~�#;'m}5��[�nL�*�Gj�(��a{��(<-P�U-��@$l,�#@�nA�e�G=����fb���@P3���.����}�ubU���\Cv�K"�@+���u�V�g�x['BoOoH!пޮ}��q���=��7.#h�DzM.��۞ݻm�7>s��.:���\qWv�l���,���-�qvm6���ء��M�tG6�P�7&��ʘNpC$,IՑn;d��z�NOaݻPp�V`�쁍�8Ϯ�r6ɜ[��vE�>cs��	��ǰv�8��v}���KQ��c������d��<���۞�m/��N����' �"���FFJ�[�ƍS֐WN��܈��"N�Wc�ۉ-�=�e�wT ��;a��g ��Wl�=�'+���1����K����oZB��w�2�頉N�Ii�)�m��	Y����,(y�ץ���N�fRagn��.(�/,�NyI�'lQ(�l{k羟tο-i�%������
z��G0�>VlV��	5��Vgj��32"	yC���U�Ks9�%�>���-,�a��f@�To*���]�X|yi�����9`��(��W�$��������q�)�W*����5��d��2�2����))0�7��!(N�Q.�e����њV�x_s$�%�	�{��KIz�+�;�M��X�6��6篆T19jc� U�%���]�Ӽä�����4&��)������wG����o�=`Cd�&y֖>���u�q����^��ŏ��^�23qf�t�Q\I��k=�I򰕦;j��g\�os�8��<M�ؚ�ɜ�lI�w��,�1�.�9T�l*|�f�\8ƈ}º���B绡4���I쪆���)t�,��:&!F�#�}��6�H�a-�{�\[;��'w��oh�Ԡ������k� �~��8��T!�f�yF�Y� ���3f�w!�Ϙ��)0�>��M��P�Ӻ�J����3��i�k_�����o���*��D�%?��)i	G�4�(�d&e�����OF��xVx�jL5�B�fG�^f"i�s93:K�/��_\�%f���iB���3^���2a%#-/��;���]�N���$*e�K֒xVNmj���fgd�&��7�`���, �E>��XP���^������۵�C���φ˅�z<���^�>-k9�탵�Ċ��֒�I6�J�s��U13$��LW-(��⒃ŏ������Ѻ��bFfK�0^7g����{3W��nR:
�	�k緎w����2t�*4�V�\W%g�/���afT�k�\��� fRa���!�S.<�<K̽.(�.��U����Vi{�6��R8H�8eTq��p��Ӏ͆�3�q+t�	�'j����s�5�Mp�����@�{��/����,�����.LB/A��#���Q�&D�d)v���h9�08~{x�ė�F��}��_w=# DL@ya��]O^��B���b�"(�� �� ��W[��J3&�F([��]\�y&!��LDJ�(nI;�d�7�� ZQ=;�$�635�a&Ʉ��B19ܫI0Vdk9ȅ�#�;�D�h���+G��d�̤f���n҅�޹�(J��n����(��iR�;�8�m�E��J[��v7g��E�!��[��s�|��V)$�2�;,,m�ć�9��zZQ�[9�V�xVNNi\��@IZx��Q�PE�`%D��UMU6a"�N�y.I�2�@�^;���Ť��=%�=�yXjI�-/�i�9�I sN6X<���{��D��ћoZ+�t�d�`���Sp�)��=iBVFbN�<<J�$Y��ͨ`I���t��IA��f��-,�-��U�O�nw�-:w�/Wo����E�4� ��tE�Ą�=w3>�U�Ǚ���񬵕�5��CKno��~=N٬~�xĬ2_j���N�j7n��N��J�c�kmf������<b�o۩�`�ۡ�Q����ӎ�Q�d87r��,���Ι/u&U�d���>G��f���
�#}V�P�C-q���\����<,��$͝]ⴱ)=��=ab̽�JOrj^�_s� ��0�,W3�nw�}�����i{Xn��hVآQ�*z�
K**�KmkHϾj���M������V=�Y��ѻ�։a#�6޿0̔��f1��}��+�|��겅"��V�%fO�Ua̐�*���s�o=-(�-��zә0�I�/��qyNiڙ�0�K����vg�o�em6rL�I��-0Q^+K����3����g��4��p�C�2N�5������D�1�V�x_ۭ��,92��������Efn)��"��E
�3\q��\�gL�Ɨ�֔L���ʸ�ic���)(<H�{5�iE�>�s�:ڎ��-�� d̯���{A���9kc��W*&�|�p<���ݍi�k'�i����!�0/�Nm�.^tڶD��©��뱴�s���c-fǵ��x���U!��9��v�k;������X��ս�83��Omm���k���Yyu����3��7M�|	�F�ɽ�m���N'���z�^��2I^|.����;O���W#���F��F��nk��=�������Yw<r][�@�_ۺ>�`�	�=�w��Ӈ��l�;�x�:M$�Z��c��m�P�9-�)����uY�~��-�F�ŷ8�p^�A�,2ԇwb�n��n�e�ۚD���~X������d��$w}o�m��	{]"9�w�s��μ��s���z��d�=Y�;�������>���7li���,�Y��oX%�����I�7k�_��|0$ͥ�X���V%f��k˹E,(9T�.q�q��ך�����afv��.(�.��+���ߦ�䙤��^>.�2y["��рL�_<(}��l��sZQ��L�&_YܫI�Lgk�I�jՔ�5<�$;��x���̓�I����W`��޸���6sUxPx��̼.����I�ߏ+��;j��QD �o_>�v֐,+�I�%�&��R���N��XI�[1�W�<+9��x�I�' "~w[n���y�k����kq��mv�����;�uۏ�-u=%~�媯�����`,���>oU�`��C�n�`�,˭���
�Ip�_9ܫ��v�B��0�D�/��N�1����펏�Y���h������h݈����9>����\�F'���~�
T�����3�z26��ȁ|�Ϭ�����랗�fB������W`la�H̃-���X�'��[��
��6��Ǥ��k/p�M��I%�voy��G�|7�Q�$��T�U�[���0@���Zl�,��tV	af��L�35AX�}���H�t�29SN�Q��}ժ�P����Ea'3!3-,z�⒃
3�nii&	m����`�%�ͺ����Ƶ����qZ%�ޫ��Y��ݦ��9&f�n��MqbV}���r	g�b �y�XP�������G3!�U9��k�>3��iG�F�f��XQ�7I����u��i��M[b�0u�XeK��g����<��Y9�[cNU�����k��� +Eltw��A��}����+77~���o�&�ŧ�F�M%&wR�Jv�eb�YI���4�^��}��ִ>�KJ3�nk�[�M�2C3)4�T�M�R�	�qǙ��Ĭ�߸S2C6ci���b4���z*�h���Ǫ�ˬV�q��w��s��m�;���Y��;<�����|<^C��t��2����r*1m������ڙ�0;�͊��s���Ó��vxbbdA��>U��A��d����������'wF�¨���tи��N�|/�8��+C	C�Ǟb��yK�U��[�:n���hT�G�P�[j���[+�sYB��b�c��cKw�B�賦���y�z2���Z�F��?{.�<�&%��xo�?��K��b���T���AY� ���6PΫ9<ϻ��G�ܖ�^~#�E��ݛݑ���䞫�\Z����;"'$тi���X���t�'��e����^�Z58H���r�����~�|{B�i"t�F��̜��{�T����GO��͋ �\5��fk?�����c1o.��8�o%�]t*(c�٫Yq���<-���1|���!���=��`xE��ϐ���1gm��;<��s�S�F*j��v��C	�5�4��_<ȳ\/2�WgS���X\N[�b �;����'�����]ŝ7�޿���x��ض���d��/������]�&t��H���{�b$-/jb��wovΦe�X���QMBn�m�����ܣ_�rn��{1����v3�f�OxÇ�f	���5�4a*�M���:Fe��H^�~�:�Z���&K8��;C�Eч��ui��8�'L,��f6-H�3e�vZ�ꥧ8B�輠f����؇��It�#++E��w2*�fJ�Ս^�Bz5��^��17�����ފ����u�O����1�Cq�_<7��冞�{�6��F��K�i�a�X�|�؇�����b�7�/SW��b���#�b2�4A��Qm�pr��/K�����$�I��E�_��(�3��sR/����4�/�ݕB���~��^����r��� ������_*3��[�xM�zO�o���fs]��Cw�����iӐ�K�(�zs�۹�U<��7]���=;6q'1p�OG�y��5ڲ�t�J�(�-/tH{o��Tz\G��b����4t��{�9���Z==ve-M��Yw��T>�o�zK��T�ؐ�����b�o\�=U��;|����D�y(�<'�G�W����M~�cn��e�Q.�8y?eBY��9ݘ�k3a���Dc��9'�}��Ԗ�0"�)��عe�=1�#���=��{^��/^+!fyO_z�����y�yyV�ƨ�S�7�^[R�-B�WvA0�<��
���9��A��4�ؘoޓ���z���k�^��FBI�d܄7Z���i��N�Um�W}�.�z1 B��w���yv�<Xj�c\��D���S�9;aU� �Qǆ����y 1�-]�瀷c��ǻ���3ǵ�|q��v�_�4-}�����}h3sm��{m�>'�^�=�=҂@�0��-�$9����,#�萌Nd��2���I�đ��#����"^��F<ػ�>�I���{����n����c���m�R��k���yn�X�7ڭӹ�ݘ�����cK��l�A�ngb��ߚ׆UQ+e\��,����[i\��L�q�9W^�������/C�F��;�I���N�^�<<��z�q����+K<+%{a�IhuH�/X%���ɗ���U����l�E���,nfa2q3Q���$ZP�O��("J�"&i)<P���KH0nL�ɖ��Mq
Ύ��,$�ڹ�(���<��Q;T(«���R���L���n[Zj8M�t`���)PUϒ�洞|����E$L"&a�m�sJ���ibVd�uV,,y�4�L��8�I���󷢗�0KS�*	q8I2LL����YZ��$�3->:���X�YԖaB�mj�93	ę�d	|d�~��DD� <L֒-(��餤�C�3b��s3�3d	s���`����X%��b\����B	X��X��-M$�d	 F�u6�iB�ι�(J̝�T�!��}��81Q#��'���'"��B$׬�wM�5�ˬ��J���5�]s�ǵ|GIs8��seXdOO:f\��gf� (��N����Y�T����Y!+��a����$�˺��Ff�ϼG����wo%�2೦�1[��{m�|� �:|;Nl[�_I;M���ٟ��6>&a ���?2�8p�)3KH0Kgv���¾I��j���->:g��,�e΍��P�&�8���H��?�����������niax�;{n��-�⻈��w{��k�､]�[[w��BVg~~|V�,(��٤��G�3f��L��D�縮 �Q�'��"@S!�DLIX%��ͫ����_� Ix������JF_MiBTd��֜ɆM����:G$��Mԣ����Q�㝙�KI0Kgg^���!�fK�{;�|%��t�������kY����)�&����I׆Ih��}�u���+7{~��E�{4��92R2H,ͽ��=���&��"$���:��<��U�X_3'd�I�u�Eh�ݾ��L(O��U�	Q��n/�{uȎ��}��$�s�Dl;T���irL�OQ���vb4;�f7AY�P�������=p�8r�3��>���	���z,Ջ�Q���U2�Kc*�����q��q����kq� n$�֣k-Z�ƨ�eC۷#�n�X�Cnˍs����;`8�c��⊣��w���m���� c9�������c�n�Ln����s�Y���e�n�� L:���Ҝ��kgq$���]�C͗W�ĸ������p�ܜ��i�ʶ&����Lx�r�Tm�(I,���U����Ⱥ���jl7�i	�佮���Z��8�ۍ��a�d��+�����'�
�l��[Uw1N�
!���ni�J��/o=�\MŴ򫹫/	X��ۮ�Ǭ�ׯfma;H�5"4�V4�ޒ���55>n+mreJ�Qٝ�4:l�>��,�zwJ�L�5��������xKO��wr�Z�,Jx�z�������rI:K��O��ur�%f�^�a���K���5Y٠s
A�O0�%�b�h�Ln���[�V�2�q0%�����`���鰣
�7�غ� �V��o����ձ%���Ⅷ��s�II���n�, ÒC$�f���\Y��jvt�2
""DĽh���W���I!%29�zH4�gO|V�%'ٻ�XX���lԻ��[�������hͧ��뜅�v6�x8�g:��I�mUA:ϖ��Z�y50���-c��RRaF��E-$�-��+<+''uW&a&Z%�����I�ӫ��\w
D�(�)�3E�"6��v�ʸ�q���K�	0�u���/*�F��4*b�	F��l!0��q}��Q��W���m�����\K�a��~T�eeg:��]����� Ml��#��N)ɭ������y����{'��߹��8e~/ĥ�s���6��Ec��xy]��Zh�8e��
{3nia̘I+4Kj~��,���%af
��U�XQ;�xQ��ٛޤ��I�{�iBVzwt�5�&B)[�Y�Z絥4�ִ�2��E%v�tR�LٍҰ��3,vd�>w_��KO�h%<��d��w���Y�̽��L(�f2���\P�9�5���m����g$а�?/�G�nx�3Ps.�NE:�lB��;�����q�.�pr��������ߟ����r�34���,~�U��
���+D����ҹ$��`^m�H����P����Q�@pq��:�i����:��2�3xZ|tWy�(0�rs��`��n��30̨I/��'w�~x�N�Ǚ
Ei�U��,���י�J��G}b����#!v��.,���ˉ˄(Z�8:(M�/]�@� ���(;�M��T�⻕j�jX��Tz�..��т=��u}��P��tZG�j���8s��Uc�^�ɘ���i�
�Q���tB�!�K������3&��r�V�%G�s^��ac琘aL���$���3;3*;����%�Y�Y�u��KL�I���y��������Im��9C�
�wⴱ)��P2K��ⴱiC�o����������2ޗ{P�;�k��e��nz�k�w[��X퇧�\�8��D9���KK%Yt�x�5"�IG�p`����X%�Ƿj޼+<Q�{t��	���>�w*����#����/������$XY���ܙ��J�(��祤%ӛEx�³jsJÒa3'->3hB��L��rI��z�A���d��A�
}�������7����^9�}�o;Ǌ��ࣣ�6"����ɐ�	&��� �Y=�ʰK:��V�gN��E�e7+7rv�L�1Iٮ��v$�3�s^[�ELO�(QP#�d#D����F,�9{P6�����ϴl d=��n7�:g�Gp�A"��j�0mkuD`3-A����i�515�j(�,y�1J�d��	�8��S��JD����M��X�$������V�G�x���g;s�k��kJi�fH�J���M��)a	l��XA��~I{��m��9#�Ste�-(r$s�[v�Oo5�<;c����J[��L��1��浤�zF,���R�i��Y�K����Ϯm���ї:6aB���W�L$�	Q���5׎~��j֝�`@��{a���K93;3h�P�F�tV`�ޝ���Onսx\�%'�V�C���V�XKC5�__�M纳oX�s������i��))0�z{JXA�Vq>��b�i��mm�o�Zi%��߻�W�ZY�;q^�(�ؽv��9&,+�w��Ĥ�P�҉���y�ILL������E%�9�	%���KI4J6;������ͷ���z=�-�_��Tw�9[c���W��IZ�)���q�K�'\#1�v�E�<T��T ��/$R��r]P�x�z����߿{>�v=��'c@�C�)L�;F����e�h�Wko)�k]�t>ܕm��Վ)q����z��`p���x�,��wh1O��c�2��cN(�2��M�h��=�n<ݵ�7gn�V��x����lH$m���6� #�+�kQY�H�0Z�nF� �r���tl�{�z�9��-�Ԇ���3��h���MMO���LN�D&��f4
[-�����G�	�W�Nщ�L����"Ɖ}u��b�	���C��K��/a�Ö��y ��7`�6S�`o{���R_&�bE1�h����{{�lb� �fa�ݽ-P�&�%CV��-e�j�Q�%DIFQS2��Ǝ�u׸�͑O�iBTd��_��N��eŋJ+{�IQ�?�zg]�lSRYe���_]8ug9�t�"J���u��->;f�+��[��s3	7�f�O�k�&ߔ(��"$�,JO��Uab���͊J9�;&l>7gz)q&�F�lVx_��~;Gi�is�U�]kQ�hz������(޽�m ���^(nfd-*�K����g��_�!>�Y����3*��ř���i�0̜L���� �|mwYX%���[5�A�fż~��{QI�ca[�aC�9�\���j��us�:��
��$�~{�����a{D<<���P�Y�:{ⴱ)7k5V,(ݽ��d��L�2Ta�]�KJ4KܾFȠI�j��m~{�w�:��bOó�%�Ǖ[=Ե��d
}
6�։�"�[�{�IF�
o���"1�us�ic�09����r*]�+D5[�x����L�]�|�
��W�պ-��5��$|.C_���\�����qr��.[��׌!�+Ll�S�(4#�R��.>��fM.�i�gJ77�Ҍ(O�z�̘L�Ĭ��n���KA��_�|>�x�=�|���i$�d�f�)��+I0_]�V	af�:�N�H���+ܓ;%c&A��ÚP�����I��٬(Xs26���ⷢ��7�N� x-�*���|i^^��{k���\���MX��gOY^�(�o�M��c^ֵ�f��o��MZ����*#��&\=���J�[���'3NWu�I��w�{���r��I,�U�%Fw_Mid��IQ�n��|�̝2n(�(����m�|��(hQ�Rfޗϗ|F�t�eC/	+��y:7ib�N�V�%'۷���I	3|-,zY���� ��J"T̪h���K >��Q����C���4����Fp���^�A V�ɞ�br��� d@b9�QHa1��Ū�ie��4�k:�P[p/��b܎����ݿ�����[¼W^����ܶnry}�(C�{�h�N�x����m�ز#r�L��jj���'~��!Y�+p�Mr�!4v��P22��0L��6g3$�	��S��z��*7��� XQ���JO̄��ͮ�]}il��ѫ8��q�m|Nf��	a�$��#$���k&<�O��X��z�K��n��G)q�iχ�sy,u���N�qGe���W��ۈ��9��ۇe�}�i��Z� F��5�S�4�,̜إ��%��\�	��L��5�ZY�<��be��R��3���[[M���&�O���\V%fϳ��E���_:��2�Q���c�����-]u��}{לu�̭z���C$�xޞ�kE&z�:���gc�.$ǒR�az"B�"����&eGWo*���S�4�,̜إ��}�w�>Ǆ�\�׻��j�����{����(X0����9I{�
k����7��Ox����������gX/cā���Ԇn7D'�q<�����s�˟�=]f�QF'�9��-坳��RP����F�}u�V2[���v��Y�M�l.����G��41�Q�u�@\� ��L"��dp�usׅ�93̶����4�>o|�℥��:�k���p��*s��c�jث��v�+�G3����w"O>�á�;���k�=�G��XGB�,Bt*ć�>t�\a�Q�:�	</�ݯ�����2Z%��]���ǫP���]8�d	�"*���>�oU{���7�Tw^� ZP�Y�IA��͊Zs!�	h�c�f���U"���2IC:Ƕ�g�ߞu�����i^�L�2��7�n,����%�����A��2�8�{KQk^;z���I��ʖ`�>9$&�L�ow���{�Z�"B&fQ�I⌇��lI!$�d!���ZX���}5�
+6)(<Q�j��x"���v��`<�!�t-T�!b2���M;ى��΍��՛�{��N��r�}5v������N�l>��8Ի�g�@�:1���;���(��o�lZ;mf�+q�x��D�y~{��{�ݬi��������;�ѥys�/0�g[�����7lڸ��3b���H_0���} �ɉ����S�Q����>wI�E[���ۏ���t(��j���h�z�#0^�n��/�Z�	�8_g��~=<V�N��n�:Ag�"���4%�d����9gO+�e��#n	�j2M��*�IT.��,pD�t:N:�DE�C�Z�v̸g0����F%
�D��˕W�̍��Q��;�P�^�1�)ODд�jq�R�p�5���z.��
qЦ��5�it�:WU+ǣ�j*�;�9o/rtj��t��0S�I<V��[5�7��TS�Z3�/N���6�-v"q6�*˕��U�w��s9�����<I�ev�\jQ��4�A��NE:i����d�u"��tPBpp[��%n�Y{Co��!U[��숩+3k�����m)����؋��=�Av��,�{	�z����ٌ��4�'XUb��ɮ����"���*��TU�2�Ž ��f��Q�1U���RV5Qg7wgy�\���ci�su�Uܐd\#�}a���WH�OF��ۜ����V�zeomeՖN!^�=轻p��t�]��Za�*��gtC���=yPs�"�umZ�Ί5��r��#o��͋�'t3�L��i���>�#����G���b��g�';=�뙹c��B)DDq�����7q�B����j������]�������$g��d+����/\�^,6��h���N�v�ͧ�ώ�/k�]�n��۞c�-�xy�v�����Ǘ���mt^-v1=��6��1�6�7 �lt;*� �\Hp�E��E�㣌��J����*�q�!���� �Ɏ�3�������u���X-��v�zqŻz.\�W�Z�#���`wGΝ���s���	���b�wm���0@�ֳ픇����݇rvų�[n(0�=���G�k]k��ncg����\mfZǝ���۴��8��"�7E�wn#l��u����g���7`H.�n�l�y�ɝ��G��[��ܷj�����u�\QI=��7Cג띲ö�%��m�c[�n۷<ګ(뵬n��(��� �I�Fy�nM1�rks���Ο<��{Yݎ�te��nv��mΝ1�Ҝ��3z��di�����y��vV�Ӥ�q�8�Ӟ8�c�dє�s�ۯ�8!��XBH��~����$^�����9��89�7]zn��.�u�m�e ��nݘ5��s�mɍ�1�s�1����rts�\�=k�q����Gd�!k���S��Ȑ<�mʙK�����7�]�(9K���tWp����i�3v�*�:�}o�����\;����G�;C���s�&����e]�v�n�D���^
26�q�xW�����K%Ѫ��Ruv�͎�^�n8T���j�N܊`�էa��^�;f�\�φ��i�F��]�4<\�-�� br��xR�i������Jq�2nH��x�W1d�gu�m��q�un!��0g��磏l����Ka5=��e=�ޭ�Ÿ�۱۔Q�ݐ�-"��$�Fu�t��+��=xU:3
���k���������'��-��P(��A[�x���p�m��vd���7��i����n�E�3����Jn۞��{J�&N:VVV�z���x�ju�d�6���ⷂi��͆6��������֤_/������kp�}��ճ�N���{�CSW�0Km�,w0ч�wv�;˷�}�g��t�o�l�Z\�A}�I~���C&,�Ù�껵&=���5��z�k�$��]�zw���j��!}��hM����zn�]�D\ﷷ��R/xӗ��p�#���7o��}��;+���Jg2�Q�2z�cUf�6�?-9�Pcr�\ė7�f
;G���8���|�e����%�N_��w��=w�<���9χ��v[��xt�M��V��5�����'�-��wB=�q�u�������.��-��6��G��8N^���.]&mK|�\���c��AG&yo)�]L=O\^xA����IB�4eJ3��k��˗�8ͳ���6�NлȂ4,���G�)������c��aY����c��7w�4�{��yo�m��m����u��z��7�ty��;�uZ{=�:���SBf�Ə,��_{+��l�-�ȫ;����)��P$KPO��S���xʹ�>�f�A��w5l�Kov�2b�m�d����q��6�}��;0��Q�t��3���9�8��ke:˔�`=�u�0}�pcS+)��H5�[Eީc0=���/{���K��<����$ۏ6�}�a�8��9�w���g3��)������[A������y�{=�f�m�K�򛵳�gM�����tw���:AҶ==�u*��oø�ĺp������Y ��Þ�oW'�kt�����cvԜ;��0���v�M�=hٲ82W40�8��ۗ�X��枫jDDhHU	[D��Ԯ��b�+-;Y��\�lpخ����^����]�Wyg�&rz^n�#�͋!MA�gw&O!���y�I�s[x�Nܘ�t�g�v�\vwb܃�Σ��=��1�cq�%��)��N�ʜh"��+GH|�?��;��+a�eF�<K*��z�τW����}�@KZ���	7�|=�{o��s{h�]��&���s_�Y#7�=��}cu��k%4�5jlY+anW{������h'�]�û���~~}t����Di�qq��K��L�����:�D���Ni_�fC2��`�0�k���w��G�8�����+l��cHw���ZrHI5�O�^�II���ۚXI�^��+�3!H� M��kH�$p�Ҫ���]c��j��|ç^�9̗̐��(����I��ʴ�ac��ucq�VB���%^���֗����R�M�$���X%�3!2[|;��q��̻rz��m���Z�
m���׊�dΠ@�2m�����igv�Ω)<H���K	0K��ɽ~�u�Q�\A�',ᮻgD���H�2������S"�"%�!��X�e���!�31����da�?b� 3'�k�2�FT��2&�M>t��ibRyO�o�$Q��)
�Z���9ۚέ�&W���S��=�Н����s�=Y�n��Ǻ��pk�!c�WGA�S��^E��U�FUj�[��4�F���gN�Os���\�qY�r�u��b/ɛ�q�Լ�U�G��ُfo�iYp}!ѝZ�lQg�G'^:���\�g1����i0��K�Ó#?�ϰZ%$�{齊ZI�[�����Z����kZ�^��'�)H" L�Y�][M��X�����d�'2o������ign��RRx�����j���w"bU,$�L�8�Y]�W`�'gx���vkb�Px�d��ڎ�mq��k�<��eW�����x����j� X}���IV��RPafFoM-(�-�ۊ�O
�`d����w����N��Ţ0Z��$m��]��\��=���4��X�/����K�Z�4�}B�+*�%���_�"w���fm��h�/f��\�BeoK�4���|gX�_�8�Oą��Q)�"EI9�L�n�Y�3�KD�q,��U��/���z�,,͚٬&a`�*���x�܆�(x����m,��O��V�%g�[�XY+�6��y����&�����YV�6��3�g�
�Nl�Iܬ$gZɁ�#��K���^��Оn&�x�R��z�����3�L��J����嶹��7��_z��q�$d����=L�Y�!a�$�\�AL�8�����y�!+�
����=�4{�oM�KDO�Y��n�G���hq�����-����α��I4��y޾U�Z|zgx�
��[M��s3�	��~�|���Q�V
ۢS��#���$XY���*JOrL*�-��T���,��z���s+^�K�L�(g���� �n�Pa���Mn�{��{9��p	����=j�{Q������|�'��O�6#[V�(���0�^�ߊ�Ĥ��vk�B�%b\xZIU;�IA���h���UF�X���z}s�֔ZK����W/^�����d�ns8�	�^���b�h�Z�*t�����������\-�d��|2�מ屾��r��F��d���+��I���Z�үZ��}�;8Y���o.�ճ�y�]
K�������!D3�5�B�*��N�۝C(�åVG��G^���t��n6��)u^,ܺ��(ỉ�e̚�0�a�<�k�fJ��6�7*~[��^ҿv�ǻ*�`����15=��緞��{a��m�-���n�|���T9�a1������Ɋ[T�S���>�͝�����P))^��bfzv�O�&���Õw�י�x��xl���o�-kʬo�wL**	p�s��կq]t�;r�\nz:��u&�ҙ툒y-,.(�6&����3ӧ;����Y����r�����}�@�Z����vRF*WE\۔|��yó~K^֖��辝|���Տ�zcug2lfK� �:�����0$(�;�6x鿹����$�����㳇�s�}�i���q�$x���?��bI/�o����:��}Y>�\����:�K~�ۋ��ޫϴ��Y�Jd9ob{�������]��}}����Jo����,˕R�߁R5ɛ�����W�.����`��.��Q�dB��>Z����UD����
��}�k+.m&Ն�A��� `Ĳ�������1�\J֧;u�zCaj��c[D/��ې{n<���i�k�M
�gp�(�%�����y�d$Ǵ��7��;��r�niXa�Ϟ�J�0�y�f�/���r��b�!�۷.����q���ݻW��;�t�n؈��ON�L����wހx>�=�Q��^M6�u� �g�
�m���sm�vzw��`}W<�no�/�d��|�N���ǀ���3֎Od���Ama��m�p1kO|��d`��U��OZq��r��u3J03ZȽU9Si�\�rv� `#,ѻ����$y4����R�c�:�nq�(�v� �v��:�Wqխn���I@Q��`F����c�������/�xo��~��:���[G�,���`� r����y���imk�3*�7���{6m�}9>�Y�%�KHM�/��O/�U�=����U�����.[;=�g����Wt�gg|����	�`Dj�j)i�Ϲ�i	i~���/g�w�u���;;^�M	�}���Ѿ�uó�91d���9����W;��KWKT�99��]��>ݺ}�W2K��#�CH�P�R�)F�+�]���<�{WE��&�x�w.�G������V}�Pt��p��߼l�]���6�'3ӻG32�6}�7z���� 9�B�� ��gy��{�~��d�~ݴ�E����&>駤��g�z)GT�'�zkP6dCIu�g��Vl�f���
�*5>$3sٕ�V튃9i�F����{�ۺ}x&	þy�����&Z��B��4���zyn�b�:)�Q�<�C2}8�����}�.��������p�Go����O�!�� )����<r�6w�s�֛֓}/�ϑ���[��a��j�"	����W��I*��屵�8���f�l�2[���2�ϙϪ�u=j������y;�[��d�&g+c������mz�k5rp�J����8�a*�V�Fރ��ι6��-B������av{�����/��l���"��R�"����.M�.����uO�/iiu�n���������!K	���=�g��bIY[Yܺ6�#��ǯ����$��Q�/ݏ�ޟV�(8�r�:w�鵼�W-�����*��L��L9�QD��8�"b�2�N �B��6#�3�`P&yAz�8l�E$q-4}�(�`X�!����fvy�{�C��0����; ֈ�u+��B��%�-����]�c�l�yV�� KF�с�˰v�ޑj����QzQ��~��������[)��X�23!�����������O&���9߀���I/���p����?<b�֘X��M[O��ru��=���isr���t���p�7��K����[�(�j8ISr���Խv.�[�����Ѻ��*�&!�A��Kf��Jѧ-XA�PRJc�1r�屶��O���ls3|���^�O|���<��/ D	L��'kmw>�o������'{����?��`�����&DB`J��ޒ��5m>�]���!�#��+���������r��'A�DV�]��x���:{W'�ն����ಮg.Y9�$��	!Y�j'cP�=�}��lR��_��k@.�=�_��u�#G�C�^1(f�F�B�xk%��c��������F/Ͽ�;4���l
��hHV�8\�4�NѪfi�^xl�^�_���'��r[P���~��c"s}����Ȉ����_X�����\"�b HI$�R���{=<6����������c�������lm��nu��Jʦ��Z����4[�l�,vk8}s��!��S���·B���)�+"(�\i�N�vegu��r����z��n�2�������n,,��rS.LJ�ˌ�>�̘fq��ۛ��9��O�26�9�s'm����<��H����/g�;��Ϸ���I�����oܶ6a��[�db�Bb�#P����UzJ��|z�s7�<or��u��ɛ/G_u��G
7LD�B�S$	���}������洺���M��<��-��KV�a���ߔ�3��O��"�]{����K���_	����}�E��t��bPm$Ip�= �E�y(\�LǴΠ�
��|��/�����*k�n�,[j��:^v�4г�朹"�v|s�sӬ�c���%c)��7��qv�^2à݃�Ɏ[]V���8���k�f�X�Z��m=Gk<u���P�۰a�;�^Dr�r(]u��m�sӇ��u��ύ�'M�+�C�.6$��x����s�ssuw8��|���S,�6�`v�9���%ƞ��l�pé-N��tAV�L�
mM|���˪u�@�`H�*�ss%8�q���	� �>��㣃��t�C����k�E�=�y�v��Ͽ/�2-�Q~���+��U$ ����Z�g&��7N���J����n%�x4��:������?�t��*%��7˝��;ۜ����WQ�<��<��.����)(���aJ������{�`xv��ʇ.����ۖFf��&^�&�x�s��)�y�y�%;���ϳ۷Q���e���$��-�����û����/;pq�Jݍ����s3y&�g_F��wElc�~ݛ՗��K$����ϙ�/<�g�-*���G`>^.����$�*6������=<���n�Ϸ'��i^����	+�tu�E!Upi�m��1��[�M�B��ٍ�K
��Q�Z�h��Y�5LN2R�	� �����96o��9w��qw�_�0��z��FK��\?�$B�T�zbd9m>�[��+�����3�Xs�a�KnxgR�N�<��=�}6����np17|dF�+nP��C3���ݛ�],��+/w4Q'] >O���&�Wx*�)�쒀{��A/��ͱ�v��ۚ&���i�]Z��]��90z�`���5r#�Ͻ�#��k���W-�9�;��i%Kmh���b�Slt@J�$������Ց������;2Pgݛ=<o~����Î�WP�1A�[(o����I5�n��z�����7v�cܒ$�*ܾ�ӵ��8�=�� �D�A&ǥ�u���{�{�4���T�<�U�cg����>��Y��Gm�=�Cm�����q5�i�w�wn)�΋�%?~��������I�$J�4:�_�?���|r�����e9�ޞ��,�T9$)��D�ƿ��[S�f\�o��s��՛���[G}�.iL�4�y{�����J��˨���峏��W%7V����kVw[��F�c/vb��98n��̇Ǔ�2I�۪��5�3���t�)j��{79T'use��'���O�l�,��4��x�Z�A�m�Ĵ�2�oY�1#�t��ۋ!���L5�sa�)(�u�p4ܜ��2��n�N5�ݧ:Dɸp*te�
&�2�o]�ڍW��^�I�Q3���g=�Ƿ�]<�b�N���	�X��W�Jt�1��=��5��W�':�]�++%�`�%$�B��˜��{�3&�í����T�I�r&�saNT+��sӘ����P"x�N(`�jz�g7�����:@=o���5a/=����w��U�3��I}S�X�dd�*SMB[3��k�36$ݘ<�N�KZQ���uOP;x��k�eM���(�s�y�l>�m�h�}u���YBВ��y>�-��{�m)>w{�^n��"��]�Ⱆ�j��Y�	¡����L������Z+��3�m�I���*�q�(8N��Q�6�]�M~f�2��n\s���O&��}WƏa�Y	�x�]����Ȏ�\��w���%�%um8�z$�"F�^)�������s7����j�޸;2�_�d�ni�F+�s�,;�i1�����x&���gOko7~}�w�I;`�|q�KM�
��I҆�����	��w|��!�5�{_Y�Ŏ��ջS4�F�Ř�蝦pGRS6�Ӱۡ����̭=���w�g;y�}}���R��o��R�`�\Qcno�"�e�Y��V�;�pIXE�5�s���?Y����q�U��C�/s��[����:��ۍ�/B�|>��KY��+	F.�]�i�ba�����z�-�lH+�''UDh�:���]I�D��~�^=��I8}��Q��Ud{�Q��^v�y��Y�-D��J���8h�#�Y>�K,t�U=��������+���z͛��h��Z�{C9t�����C�y�]�<�o>�zx�@�{;*�!e���N#\\wۻ�r�o!�f�R>^��X�fE�I��и��[y{{����J�Gd,���/��t��x�pSÏ.��h����[w�Z6�c}��8���S����w�qH��CKa��R���Hr�sLD䕁��3�aQ�vz?l�3��b7��y��
%5�ܖ���=�䶮f�������=&�y���|w���t��ԟ�Ky�1��Ռ��tnp�7^[�O=��KQ�|�����njm�n�	�h�sK����s���{<�3�Ηr��\�3]5iė�P�	�0y�^Yj�{����|zБ]�ۄi	i`�z}�Ojpoz�+p�Ouی��:��v����W�'��,>��^%g�� �"b�G#ND��f�˹=�❇�wL�-:;�ǖ��$������hx&W�:6����7��})�����5� �r����ꣷ��X������ƾ��)p�e�Mcy0���+%k٢Ϧ�����!�4��.]�p\R�{�v���7&QGݩ]�D�U�����Y�=Pu�)yx�����{1�ܰ���֟m�:Ę��t��(~����ѓ�d*�����=F�f�'->��?mM7ܲhNGH�I��$���z}��Z������f����fX��+{��+���C��¹T9K��7��>���Kl��߻���ǝ���3r�c'�Jc;�!�\�!��x�[n3+2��vn�흳�[�]���HF�ӓkK�+��i���nA�!))����w�ˣ�͞[%���@��v���|s�u��U��#��Io������3/2Jr����_d��X��ܽ[̛̖	^�Y\��~P�LC�ND��іon�������Yz��s;6'���D�X��U���g<��$�������\}]��dth͸�p�Y&����Ɖȭu0`�t�u�c��w���.S�}N��&~�sFN�[�<X矏L��N*%��;�	ݛ9;��}�C �i��*`�+�m�������[L�9�Ώ���\LD��|-�[���p�����>�D��b��O����.؃�a/�8��]olj���U���4Y
=���w';��ZWZ���я��Eg�0�����dٷ�<q;:���-��ml㥍�����<�C��۞��m�TC���O�ֶ�ƞg�t�nP^���.[y�:mC���g�[w�}��ܳӶu��b�dD��>�9��fvL�k{���}>�|���&�y�L�f>sS��n�WU��N��|���l��j=���L��螌|���&7e���[�����ii�K=�����{�e��ߟ7VVs2Ԛ������}N.h{gQ)�)x���#7_�����Ww�\�=�t�v�w�;��:V���S��wi�Q�Ee\�~�荅�xr:�b&�[ �5�63���/.
��M����?��yi��F%��ܹS�x��di�YX(94_�����I�K]��\s���nyq�Pb.ܵn�s�ĳ4�o����>��綨�^�ؔ:�i9{uu���� �����ۺ�:�ms��
i�{f�K����i)�����:�XoP"쾈��îț�{J�&�K�#�l=���>6����z�gN���yk�6�y�nw����K�;O#���ە�s��v�׉��F�l��1���)0?�K��s$+�6P���%��~�P�䯥��x����k�q�����[�b�5�~�7��,��N�������ڗq&��� s���`��[�f��m�\���y�Ȧ�.4vv��6��5�'�X�AZ��쵷]&���˙ͧ�������7$�M���+��������;c����9�/:����C�����O�K��Gw�����b"�`̟@^��|����/�s����� ���}���6}Y�l���L��ɓ��f�������/���#2=����$��M�x��߻���:����C-P�������\�RIu��Ⱥ������m���=�/u�<I��,,��WY�#����[�k'.;C�+�aE��WD7_�|w�����2@�T��]��������9�9�~w�����ik�?>��~���d�M�`�Rzv��rc�}G/�EuR�>�δi�br�G��*����j��{��l�u�>fv.��u�2\]
}�.�V�$�+ê\�E�:c*V�}~Uq�����2���{b�۝۾����lg~�"��Qc��l���Awd<�EKݬvꌓrj��؅cw>}��L�d��wT������0 $�޾y��ƭ�%�������ӓg;s�c�2�Im{����屒o�g�e� .��ZW[i-��������>�͝:o��֦�[�}����<���en�����w�7�ֵ4�{�޽�=�3��g9����<��{��L҉��eT��Yqs��:0\m���Og�h.�+��n�/��{�}�3Y\pR�����}������g����ֿ&a3}��5�ӽ�B}�wqQ��8J>��O�|����f�}���6�\�^�͝Yɛ���kj ���0H""_+���c+g6�F�gG���r����'x�9�xH���r����������=!޹|xw)��/�G��ԖC3v�ګދL*�ڼ:�_e��6A�ՓL�1�Jf��
��^�㻎�mѢ�q��z=�j0,>�p!cYzB9j������5Ջj��s1
����{��1m���巍{��dTm��������]�\���p�ި��۱[s3bkz>��}�X�^�Ҋ��Q�l�y�WokZ�t��o�
�Z�����Ot�����}q_$d�����{7�鋳;�h�us�,�Ѫ睛l���ў�_��������I)d4A������>G�w.�g+r��foP���q��gj1�JdhO����|�fĚ��}��:[�R�yܫ����l�%r���r�i�������f��ls3y�m����$�����65�'��u L������%�mw.�~�������V�g�97�c3>�ʓz�F��Fϻp��1ݓ����G��$'S��|4����׀[��
�H������*�Mإ��0�_�VJL>u���ӻb��8�R��iƪ睼�ԫ�����ɍ�3�U����t�,���>�Y�t���'2��Ȼw���ii���<�]���[�I�π����eEn'iuǝN��m�쳌Ol�P�� %B�W���@]V��_��z�V���HZ�HP��k���_(��X���ߟ���f�����r�/v֯u��l�y���3�����/��tw.���;�?�w.�9�'fU�[�!�wTM��A��t�99������4����Oj�����A�p��f&3s���oF��del��|�g5y���KQ�g}�m���OJ�EjҰL�g��GKxx����t9s���<ީ��W��5G�v����^�u��k�������;�u��6����!jn9Z�D�A!ߥ�z���'�dі��a�_�����3V����#����i,e���⎮Wh3��>�e�ݎx;+�FڻZ��(g�2�����i�<\Ip8�np���V��7=�Be�"98+#q��Ϋ��I���6���N<�k�������]��\^�\b��mch�MЎx���x�9��7������W)[;vM�k��h�c(qɷ=�����s�s㷛 ������L<q��흝�{u�Ӫ�?��V)ְ,��Xr����]��x�d<�Yݷ�᪽�9Y�)�{!���rhoQ�jgl���Eb�м��t�6�u�S�����tn{;�X�x:�U�5eH	ת]U�ִU��vV�N�&kc+����ӗ�'��?|<)�}��;�NE��`YQR4�=���:|s�Is2�ms�������+g'W��c*`�տxO�9*TK��$��;�fǧϛ��̒ĴH��ގ��ܟN�B� �S�91<J�{�%���{�^��}�kgg��C�� 1��~ȹv^��/�*TAE e$�4������<�x?�ܞ��讏?�v����2�9�9�P���<A�ڮ�z��i/����I�]��k��wA���kIBc�Q�PB�����w�Zr{k�-�k�|�������<����e��r�D����W �N���N>�p��۩�V�\��=Q	�P3v��΅t�I����X�F|�.���,mqɏH��و9�w��G���G�)����y�l��SZĲL��F�u����_�;M.h��X�Jr[W��G6����=�Y<�x���ذIVt��ft�G��t�+:���ml�o��=�����|_���PF����ϻ��'kS��� {O�}����[Y8�m!��[����i!%��������}�l{�%��Vu�OG��\�ߦ$"d��D�G�wVnW3(L���md�u���nT����3gwκ�QL��r�����;l�l[�R�q�"�����8܍f�xp�$������n+dD���׽���w��O���ә%l�/<d�G{n;Gy��W%J
��Kٳ�Ý\���Z���^�c���~22M�j�L�$�(�s��&ܶ���9=�;6w�:���{��s��;�#�j'�cJ{=�fx���qz"�a�|���S�U}�,Р�WGA�熭�X�,C[ ޯ	!�B��KB�{��9��~k���X<�!8qL�u6yl�ᘓ{7�˧�*�����2�Ò�.ށ4��m�[��㵄�a��_ �Wc+�]s�O��8&
�AJ*�����._���ֻ�Hr�}�O�����NN񓗯�.V���\Jf&3s�ح�O3,MM��O�9�<��Y��<�ڸ��ϝ�Ρ�����S���σvx���c�6{^����7su<���?~�{�{��������D��	BRi9{��=M�.��e�f�̗&m7��[Y=�*Ɉt�e�@93;���S���e��v�lm�{��7�;����5֗��,�,��h�D��d��y�s�Ӻ�y��kc��u�}��<������(;"�-/=�k�Ff�{�j�$����f>m�Ϫ�Tﰥ�T_Y_Op��Y5P�1���^s�Xؓ2�W�BwS�1�b���ؾ�I�wXŔ',�g��WZ����z�E��!�]i�����07H.}f�C�Vn"�ExP�E�!�-�L4Q>ٿQ�K������;6�̕d�H�^P�#0�g��sN���{����-]&���ˌ�)�=|ɽĻ���R��
Xtg��8�V��R�v�x('�,�9x��m��3�:?���WU�լ��v����/|�o��w�|�î����{����쯗Jߧ��"!L����)L�[O������8����w9�NgM�i}�Z_��{o�d�VW$�
T��_�=��˝��?x�>�gˣ��ח�qmY�g�*��h2R���i(d�ow|���o�^���ns&vMQ9ܹy���9#g�j(2P:�9�}ë��x �ݿ��~�-d�ræ�;�� ~h���?�����չJT�����*�o���9��=�}ϓ�*�D�2�:8W=Ѥ\�%u�%s��UK��H�h�'=$.�u�T�]5%I˗���q�.�ϓ��2���JQ+5m�����O�Ǘ�ׯ������O�����]�8����q����W%�?�����z}^W{�̥J����g��>TU*�
�U�4p�g��w�:ې79�T��k�m��������)R����w������:�N|�_����y�<�^\�8|7�y�N��?����G�����W�q�����Vj�U�5���љf�efLɚ��֌��������1f��K�Y��3Q���5f�e���0��ZY��3+2��d�Lњ����4fMa����Y�Z��d�,�֌�س&e�Z�j̙�e��e�����L��Y�Z�յ3Vi�3j�Lֵf�eff՚�јfkFe�3Ka�Z՚��if�if�Va���2̳Vb�Va���ƴf��0��0̳S5k,���0֦j�՚�Z՚�Fh�5�2f3S0֙�53Va�3LљfMd�f�0֙�h��Z3Ve��SZ�,�c0�L�i��Y��f��2�5�1��3V�f��ɚ��F�5f��e��fZ�i��fј�fY�i�f3M�jֳVi�f��2�f��Xf��4��Y��kf���3,ư�f̳-e���2֙�e�5��̳Vlƶi��f�f�5f��c36cZ��f���5��f5�٬�f��f�,ִ�lf,�1��33Y���5��kY��5��̶33��5��ֳVk5�k�i��Z�5�f�3Z�k31�֘٬ƙ���k3Y�kmk6fk5�333fZ�4�f�k33��5��k5�ֳ�34��kY�5��Z�L��mfk5��Y���ml�6l��kffc6����k3Y��5����k3mcZ٦i�����kf�f�ffmm4�͛Y�f4�c3�͍��31�f��fkf�ffk3f���i��3M�6f�36l�lٳY��mk36f�͌�Y�f3Z���5�M��-���1�k6�i����Z�͛6�6��͚ٙ��͛5��4���͆͘�3mkcY�4̱�����3ff�����3�fm6ll�٘ٵ��3cfѱ������ͣlfl���fmmmM�M��3&ճc[fֱ�i�e��c4ضlڶ6���ڶk33L͖�����l��mfl�ڶm[[-�͛1�kfѳem666��f͛[[5�c5�f���m-�M��V�ڛ[Sfə�fŴ�[&��m[I���f��66��cfkf��[��ڶ�jl�ɳj��ͨ�6llV՚�j��mM�6����l6��Q����16���6�66)��cbmK136��Fձ�l�-��jlmV��mKj��a�6&ű�ڭ�4���e�ڛL��[I��f6���&�6�Uk,�b�l�[Y�1���Y�el�f�m&��1��fM�Ռm[+Z���m&͓f�5��mllf��j�ڙ����6�ձ������M��dƫe�Mj�m34�kic66���͖�ci�l�k)����lسF��8q&263)��16i��Ff�mZe5���S4�5��h��Ɠj��5Ze4f��)�mF��Z��&L�6��j���&XڛV�&�-�VSL�YmmM��jj����2��ٵ�hє�,�ML��F�LZL���ML���Vզ6[FƫI�)�ɚ�16d�b��m0�d�j56�5L�6�2���VV�ѓTɤ�Sjj2��L��SFSL���MS&�+)����cKjŪd�ن��M&�S�&�M&���SQ���je44�5L2�i42�4�5L�����&,����SSI��Ɠ&���Ŕ��j�d�5i52�4��L�M,�M,�-&,�VS��F�FSSS�U���b�0��N%��I�)�)��`���i2�YL��&FSSI��2�M,���U��2�2��LL�,��)����`�j14����MF�C)�I�T�i5MM&�)��hi4��M&�S+)��j4���,L��M&�)������0��MF���)��d�j���&���i2�L��%�����.*b�hi5LM&���I��jZMFSC)��i4�,��I�j��S��e4�MSC#)����j2�YL�&FS)��j�M&���e4�M&���he0�����)���bj�MSI��j��&S)���e22����I��j4�MSI��e04�L�����ұ12�L���)�i5L&+Tʴ�MV�)��j��V�R�h��L�U���be410���MS)��ae2�LMS)���hi2�LMS%��e5-&SR�e2�-&�)���j���)���ae4�ST�ae24�VS%���h��L-&�T��eL��#)����4�LL,�KI��4ZL�ST�iYMS*�e4�L���ʵMSE��e5L�����e24��LL�&SCI��`i5Z����e02��L���i0���&���e5VS%��i5MS)�e2�MF�R�iYM&S)��e44�MSI�e5M&�)���2���L���be5��%��i0�LV�)��iYL�S)��b���S)���i1YMK)��b���MS�+T�i1YLM&�)��5LL����e0��YM&�C)��ҵM�)���h��V��I����be0e12�4�YLM&��i1YL�I��bbj5MK)�I��`�iZ�+I�)��h��LVS��2��&&��e24��ST�aj�LM&ST�de5YL�SQ��e4���ST�eYM��E�j4�L�F�)��h����SCI���e5VSSU��e5MS)��j2��&���Եj��25�4�4�%�S2343Z�1Y���bfS4�Q��j3I�����CX�����5�����L��,��L�̍j�)��Űk+1fL�f-j34�������1f�����,�fSj������,�k+2������,՘3ikC2�I���M��Y�fdfL��3�f&if��kC53C4f�YY��3K0�Mif����)�L�̌�̭j�)���2���6�4f-hf�2�&i5�����Y�Xf�d���,��3Fř�̬�5f-hf�5Y�1kFjf,��-a�]ϧٹ\~Z��W���T���{<gw/��>Z���������s�����o���}��R�W.��r��v�>���}w���^�_�Nޛ���u}�o����������N�O���)R���mg������~:��ߋ�^����T����U���.����Us;z���86p��������R�4s�ӎ>���ڿ��;�:v��ϧl�?����qf>:�7�7�3���ȥJ��?[�}�C���^����U�w��;��×�A���v���@���<����w����v�9~?��J�_W7?K���?g�yV���U�~������|��z�;+�缺��u�9��t�K�q�t����W�n�?���x9����~M�����_����*Uy��}������n����N}�����=�_��v�����oO���|(�U�q}�/��������ʊ�W��{�>�������7N��>?7Û���_��{n���PVI��O#xg��N��������H�����      -B0 ��T
                                    8𒤊��Q*�%UB�E!TJ�P�B�UH�UJ�!T��@� ���)�I*U%UEI*�J����T)$DJ (R�*�(@��R�Q *�(���EEUP
�J�T( J�

H$)*���DE
�Ǟ��TUB%*���  �ι�������`9��f���m����o]�	�礇���B��<�P���P���[�jW�]��$�;�]�<�mF���x;#�I*�J�� ( ('��z@�A�k�� �"��x>�A�:A��N��}�: �>㠠}�AAC��w�|A�h(4|׼*��nx�@���
R�P��I�Yv�#���B�׊�@*�T�^�	E@�R�� J:�7w�S��/3ݵ�N��`��q"<Y޳���c�S�w{��(��皆��k ��nEɝ��iR��&{� ��-�՛m��T�IU@P��
�*�cP�.��p��9�T��s�֚�[�z0��j���y��`�ޞl yn$��n��5�Ï3"���郈P�L�J����EE
�*�����*�%T(�R)EQ z��᳼�B�-Э�:n��t:��.��
q��x��@ZǏw���
0�=�+�^W���3y�ZS��<���pORI"B�RIQ
����hs��w[e�����J�\q��A��*m
�X]�ǧr!�'|"_z�w��Vv8�ޔ/,+�1���ч�Wz�+Y<T�"QR��z�$��
H��U.p�Q%W8%p�u��3��n z�޻�I�k�w*�;�E���͹��U�q�e�e޷��W��i���J���T��j�XS��rT�H�R��� !�{x����޷J(�RI�;�W�;�G��/Use�6��t��A'}s��5b�z�V4���d��޷�By �B��z��T��%%ET�-�P�JTWrAn�7�U�w֥x�u�s�!N6^�Dn�*��*�qza+͠�-K�{�z��A�P�W<:
g��C��6�� �*�JUITQIv�w�S��&w��lP�=J��u@��=��`{<h,eh*�7y��s�����!/^�=OV���{��z���[�g�[|                         ��JJ����    2S�0I)T�� @h  5?F�#MR���!�d��&# hD�J�	���h@��  =F�l��H      !I4PM<�4�OI䌀=ODl����~_�$���~��������O0���8�..7�:�;�� (��qǶ��
�*���!��TO�U� K�� ����@@��������������4��*��g���
*"����O���Gw1~F "/���g�x�_�x� h��� Я����O�)�/�<J�9?��Hu�&�!$N� w#��?�P;�;�MB0 u��:�8�2��r�G�Nad��H�J���^��C�_ `B�}�M�J�@�����/0.B�G�G�^%u	��SP����4"d d'2�
D�T�	@��J�%N�N ��)�q �@�ۑ29�Ndz�|�z�PP%�`C�w*u-J'&�N�^�rD���/��w+�
P��D��@�䚐�
@�A�S�P��r"y ����܈u(�� �	�q(�=��S�C���W�)�\�܊{ �B�0y �@����^%]@�!�i�NdN�( �'��2���CpnD�����%�ԁ��]��n�M���O ]H�"�n]J��w�7
{'�P��̝B=H�+@�#�y�8��|���u s@jD��z�2�N!L�2D�}����E��CR��sI�	@�.B��%9�28��5�J��{�'R��:��J�.�H��*����0�0�
j_%W���Gp#�d'R��p'�&�N`ɨ_ R!I�!�&BH�p���N�O`J<�2p2	�ĉġ�)�#�&��a�@�'R���.�}���C�;��C$5��( {�i_a`S��Wr�̇����@�W��ܪs+��/:�܋�_ B�"4 /p�2'p�Ru�� ���aN$dR��rG��rP2S%A��U�D�T��UԢnU9�W�9�O$!y�2T7=ț��Ի�(9���N!z��MJB=B
��PJTF����=�c&�uٕ}Ig	H%2+w`�p�3��g���ga�]��)C��f*h��׈�ǎ�4'��p�+^O?i�ĸ�y�mJ֯_{�w<�;w֏�]��F�=��}'x��X|�����M�=5q��/oOrgr��?(Bŝ黼q@JP>��>��h�K6��&��\?T�e���s.Xٙ
��Qx06bH���1�.�3,��t��V�a;�����}�=�> Y	ԡ�'r�Jd�s Ҝ�=@>B�	�
d���'r%"w ����T�D�B�}�)D�!�S�D�@:���SPȜ��)��K�SR R%"w(w+�N�e;�:�9�28�:��%x�r=�=�5�	�yHjP�SR��J���(^�r�(erJ� d�"y"jP)J�N�3�_e{���8��P�C�!ĩ܀yB�J�7 d��)S�^!��
P!��rR�d�ҽ�u!�e{��:�|�5 u"u u(�@�ȅ#��� �
w �J	���� +�_��cr;���?���fA��F�	W�,\�1�{��F �6���=��J$cX��-y^�T�eFO�(,v�cڡ��;3�o�ͬ�{����u���S	�ǡ>0���Sm���m��.�w`gEޟ�:%�a��x����(3��deb�5����4���7eP��jx�z�eC����b�+��L��v�+�
�rA�Ԑ^ܝ�Xb��v\e�;(�ܰ���|��(x�~�s���L�ef��P�S�%�E��D,�53ol�����c�6������q!�d"T�3�
�x��4�Xu�ćpmDm�-������Dh�Y�����P����[]Iy��5��[E��o����=���r���m����=������o-�y�}㉼�f,5WƏ, ��x���A����N�D+<���VƵ/v�����\z��Ѯ�ɩ��Z.*ؼE�aʔ���!4Rq�������hgøzKt��0��O�8l������]3� �:d��DzŖdMޚ ъkժ2T�������Ցe���G���wVM�#�[�5Sw`ѫ/a4�[�f��L�z�釸K�;��ln�9��Kov�[ԋ��5���;���r�Oy��.����|�!�\5�6t�䵇C{�����؆�I�.���,1^�kq�Ô�0���U�2�l���v��5ܡ�H�ss�Q�f����atz:�О�]ܛ�WcNw;���^�՚�m��ю.02+;Eɽ3h��9���o�LU��v·�I��(�� -=Xvݨ�	MvԲ�Q�C�='Xx+������=lL��W/Y��gNTH��8R[J�%XM�v�ܱ�x��a$����`��xD](󺪗�s۫"i����E���J����Fs ���Bf�2p��M�w��i�V{�J�p7q\Xv.͚v�3�l%\�K�tw.�3);M���؋�MD0�`��Ŝ����N���/AЋ` Z) f�^V�j��=��r|��:h&v�&4u��~����E���/�[aZ���a}w�$u�nXlO�V%1��&$w9ö��ۿ�S��.9����!9B
B�@�S����֗f������s��SVv�k䪃@9F�B�
���8�\�]x���g>3�aB�s[�w�ہA�lDqe�M��k��u��-yJYݶ;�9����&F̠_~��
;��b)�wu� �VcYtn���#W�nǻ�{9	����q{ ㆺ�\{[5�v������O쬜�E9;��qjLb�80d�U#�$�B4�pz�,[ R���Tv(��	n����x'@���ڲY�Z��ݜ�c8�,'6��Q|wv�GNɒYd<��m�o*��U���!��X�Zh �z���ѡf�"M����4voN�=T�.G�������dՇ��ă��B6�������]ܚ����3=߻��{��Ӹ��J��S�~��c�k��q�Z��+�U����.μRvشJ�s�/�7�i!)�#k���)�OGpMG�Xs�dD��X�#�Mޜ_m�I�4"�wg[���
����mèE�L�H��:6/Kݬl��͙[�5�N'f�]�H+�`���pe���'S�	�a����r�H>Y:T��U�n��5�Y'7�2��a`��ߤ��3�c�̹k�V�r�|��ð�G�M{���5���3��y���=�f,:�Z��㇏+�^����K��q9��T�"�97�;����q8f��,�$�.��Hb�4���Sê:sv�Z���1Y5g@��uͥd�.U����u���)�׫^�ݻ�'�`�3��cw��u��mi�Vsj��b�/Uk����;Nѡu�6�$���s�>�u�����s����
'S��՝���(w@B	��;fv>B��3��d-!r�ǳO,��tK�Z���:��S� �/͞S|�v�.����㛏xdM�/c3�1@!X"��D��d�B*�$o#�Ic�a�Iv�P�ܩ��k���ĕOI�h)c���@��^���PE�N�6�F 3p�����Vt룣�7�L�a�؟�9`��nqud��qS��ܮ��3p+�.���������::^��(F�ԋж3x�g^��u=1r b a�ށ�C�v�z�:�['%cg�z�ۉ�儝�{J+�V�:���Lz�t��kA�����f�9f��TO��f�f�]3�w!\�s����lN����$��ag���f�<�rk��t�;��l�`��,i``~��J�A��]�GcĦ��5j��j�d�y3��fm=ߌGnp묂s��"b��H3�Z��s��br	�d��m���J^�v�����u���^l/n-���q��v�д�����Q�-ǫr^2Ib��:�,<T}����%-+�;^nj6[�S�(X�v���N�މ�(�\��uƖ�O6��Š��oX�M��]Uxt՚���.[��w���ɝ3n� �r]o�e|��=�1we�sv�a�%Z�{�.�D��6��q\���8�z�Z����/p��F���3��R����>ˏw�P��Rt��c7DssuˊC�f�{�����_p�(�wnQKVƮ-�E����&�(;-: �[R(��3MԺ~]�7#�Ӥ�ܸ8;j���.�{iU�`ދ�Q�B�Sٽ���a��w[�An1��&<���MG[�� 1P�OX�L�U�:�!�aA� j�6���n\��;7��o�^�.�3�@��_qh_�c����^su��a�c)\� wyG�i��g�jb�a3w�b�S� ��!�l�����~��Ď��܉�a(.J��;N큸�Ϋ�:t�sPŋ���51�������$��0,Ap+FpOCi��]���ol�y�ᔳq�\@�h�SĖ6s�p����|��7/F?Q�m<y�t����f%r]��3��{��yA�x�ˮ�l��I-��`��{7�}�V^��2�!ѷznʗ�n?�;�$��JM�ڃ��ùVv,R�:.͢��y����&�}2Q*�y�=��ș�Z܎D*�%z�;;..�U�v[�w@��c��[q��XP,.֜6Ǉh�#�wT�omՐ�{3N�^E������c�.�U�v'0@�ZG)O�HN��4%�_u�������l��G�ݚs�	��)3���HE��j��ש�έ���On���>�WM�Q�5��ԡ��TcǶ7���x4M�xh i��V;4��������'C:��H@��b�3�Q[�N4Vq@���e��jwG jt��bNZ\�w;�BҐ�8�8�ע��jF̄��cϷss���]�r�S�ް�`��?S��$7���a��
����74�UDs�,fѹ�
pMķ���Y�f�8�cxygV�csf)����?98�q^ۅ���|���{z�Kq�"��:���w7�W��[J����J�v�M��;D����X^�w�f�v�%�^vG����V1F�zx���xn�L�۽�S�`�?F6i�����&pމ�/�`8�#��7���yf 懁tW��icZ�c#8�E�x�ݐ��:�KMr�܍��N�\�rKv}�&�Lcu�ƞ��i�u]Yvp�ԣ�; ��]�S��{�>��V�8t�T��i;��2H^K�Jܓ�Ći�		Kvу`���շ{t���:�4�F]h�;�O6�F��c�ݧ;_aw��4�)��kEgh��xߡ��bmч��b;ha����s�F�����nE��R>����mx:Se@6���Nv��!�d7�	^��wm�� �1F��(.�X�7:��G����[ݑP��7����ɝb�O0�QW��r==A=����sw���b`�2m\�&�.�;�4\��f����_f�o��Gk5à66�ĳ�n	�]<Gm����&��rC#\��ڷ��P�jtfj����98��v�`��t��`S_b.׏!���>��8��+�R���IK�P�\j��.Pv��F�lT��rHE�K����G�İ�wV�~�y\}7o ���zN�sf��ú۸p��쯳ub�e��;v�ֽ ӝ������庖�������Np�����iۧH@u�ۂ�X�P�>�S�*������G{7��z@�q�	ݹ�Hn<ك�=�Lc��0!�����o�ˆL��	�� \�ǭvo�0=�v��s��Y&�y2�V#��v&�����\v�����>�:��,�0t�I9z�/����
�.�wp���8�h;�����K2��2
L6�X�C�u=��u:8�x9�%{xo@��N���3X�6�-����oH���p~S�w��A����-M��2�U���oh�K	"-�F�5#� H�hc�a�H���V�5����F��ٯm�w���pn�X��o!���մlK�Ϳ��ky��J�;�՝�6U�7s�yk�H _� Z�����P��"nRIu�{�v��rV/>�^^��[��oR��OM�$b���(i�w�k���fwigG��3���,�و���*g"���6��\츶�};���h�D����Z�h�Q`�C!lK��T�At��:�n�Q)l��7�R���պSƩ�!�z��,��k!͉{��{��on�9V���p;���w���o^;�h�V��Y�n%G���"��.չ?%U�������݋�O$p���/�vl�������±־�x��{���8�/�b>��B�C%3.��u͹�b�#���0f�E���V��T13��ʰ�[���f��7��r	���}���F�"T�>k�ʶN%	��\�wfR�h�2R�E�L��^Q�46=���C�v�uHsH���"q-FT�@e��T��0�h	=v%�]UG1�=Wd��0�|�[����s��b��"�[k�����5Z��!��O��7�V�k!�܄��
�<t��i�鈓��Ӈ�ft��.p8�.�n�i�ٻ��e���l�x������}�L8���2��7i�7j�+��q��{/+����ts��%�,�q7��y���l/0�d�kOMh�D��b �.�`�Blaō�ݝ�7 �Oww��)9m9ۡ�x�����1#���;�D�Ӱq���U�󜜵�6�uu����"���Ӭ�䃎���1>X���g)��kl���Sr7�Kk�7�{;���yo�6M����t!KhӦm�.Z@�	Z5�����Ek[�x���i�:��l��� �{p����v=�N�=ʗOTW��իH�6'�p'NiiN�:T��ڶq�4*��o^ڪy� ��ƐR��jA~��>���È麪�dZ^9����� A�]�)�or��NZI�+�ù�h���=Yw��ȴ�9 �:�rE�vI��d���N��ey���0gH�4���q�#<���7k�=9��� �0i�m@n�7;�9��:`��u�����r�8�g�nsf�%�3c��t2S���8��s��vѹ�;"���0Ӝ��;���{���5>Y�wn�����ͥ�p�՝��o]��+)z��� �0;�����Q�8�7BƶA�U溮0={�WI/	�t���u�ޜ��:i�E�t�{)
��=цP�����(R��{!,��'1�O34�(qG�#y��ju4Hῑ�Xqb��ElOsE�'>|f,��#�u>�t �f���> M�9�i�q�tlc+;n�F�#���ȴ�r~p+s��̏5���8�.���CU�R\ŪY.5K#yT%f��u���N���w>���X��w��7^�̹npR��|!��k�v��u�U�����Ƹn��Q}��ɏ$��o;�tj�\k	�l�(Ì�C��@� �,�[X5�+̛$�,�X)�(�I!)6`�zp�1R��}*����Yw�{�_;�ɜC.=C�W�%z2��	1��u��S��2�E�R��ܢ��H��U�"I�f.;C͡>�]ܶ�d�[�^6��p㗷U�N��R�ϋ=�%���md��M���*�kL��JE���;�; z��q��睝��L�w������M"��;���&3I�\ݚnM�.�ѽJ��"�o�3lI�����0n��m�j�� ��L��V�F�0�8�k{�L=y���Ju|չ<�dQbG;v.��o�y܂W�p������X.E�"=���iV�9��s��y��F�hYݹҞ��&{]��c�E���s�[4!�V6�����ݮW�QA��;�̈	M���h��xY��0Ɗ��L��\�C��;;�}��VN��� 3Y�����p'���nL	���8��iwY���2��kV1��A� ܹ�{��*f����|�0u��١p[?Q7B����#
u(�<
�t q�6��G.�م��CBGx����ǣ�^{���v�޽��	ZUy�w-ۯ3m*PEٷPU*��p���w'����`I��w)�y����!�{ ��V�@�T<���=|�h:`��ش۽b|�/qt����"�f*��K�yG*ݏj����ǻ��}�޶�k��}�r\�����7����2��^���}����z7����aӵ�f=�֨.T4ZN�'��M��I�Q�6]�Kq����xDB#��"zix���(3�5�p7OJ����}�V��`W���A�}�Vy�њ�D'���B���.v���a�NEu��fn;F0�^�r�9t=O<׻�$=W:Y�����0'ڮ��C��ּc
������}�����^�k�_w�_����-��X�sum�y����4ha��"�2�.�ie�Z�ˊ���Dp�ݝ2��-0L�%�8��݇0oLm�1�8�x�+��~��wͭyv�ۀ<r۵�Q�<�[ݻv��ܔn�N\c�h-w���x�+k�5���eLR
Mf��,k �kku��)�v*�v���9۠��:����BΡ�q��'!q��o:������찍l˴��1��j��@u�w]������i����0����%qYJ�h��į#f���T��u�����<kfyfz�5�V䵨ϙc�u$�kfӡx�o,��f�e),lf.��f\���-\�6dmt�ˢ��q��n2�SS#w3�<u\g����gn����L�WQ֭f� ��,Î:��[����t�ѕ�<�#����ͻc���Y��ijc )�6[�CF�(��\P��/��ڕkb�i�gu]�'��]�18���6�Y��F�ej�����
\����*M�(B�Ii1�ǧ�N�WU�_=�1�#:Y�T�)M5f뉣���qV���7�VB��cJ�f&aE\��h�Yq+����N��y�<��j3�vp�ëJwA]&Aﯾ~n��^�mۆS'n՛��Eذi�e���s�H$���4�qfVX!�سf;AXi[��؎zk#�lVp܀����ƴ��j�Bg^>Խ����'�Ѻ��ϑ\�D*��Bb��u�j�Z�=yt��5Z�;s�cg����ee�2�^]MHjD�	f�L#�Y,5F�p��m�Yl@���)ui-Ք��V�5�e$E��X�n�*Z�A��7j&f�����V��j�>�S�]mcO�0BC��S�67N���\�ڗ�@�[�+�S7Cke,�m<mfN�voZ���ۮkZ쮨�tuy�p�]�ʗ=��Ʉ�x��猈�����V��Jr�L�1���N�W`5uK�}�,I�Kp�TЇ]`�!,�uB3.jiA�Jj�����-fL̺.�!��fm2J��0��`6�	m�EB�x�v�ke)y��	�= �d6��z�A5ṉF��X�n�D���z�p%�t^̢�z���U�&�jXqjL֙$(��ּ(Af@�]��O:5��npH��y�ϝx�[��,�l��,n��c����ڍ,��Ps���y�5#�m�x{���OG���\�/'U��	I��u��U3. :��2� lk�,�X�ƅ�N�§nn�J����;�ܓ�=�ݸx-���P��ۘ͋$x���n�=�C����p@�7��h�-��F��*�ne���փ�r;v�z/+���!0�,�f�5��5"�[�ٸ�t<��Ʈ,ln��v�~|����'�9�����rW��k5{[�l���n� =+������UN΂w�178���o&�p���<Onҽu��t8��1K^i�WM�m�b�Aڪ�W��:]��Lٳ�V(�Ү*��6j�JB�
��1�il��{�0d�.+[Z�,�h����A���o�k>���P����6B�*����t�!
���e[�n�^m(Ւ�S��1���I��hն�ˉ�۠჌]r�c\��λB��v����{]����u���e�]�4��l�׵���k+U�k��|a(8��0G��8�vksO�"=�}��m�kٰ����㞱�KN:�[�X�Fle�6�s���9�m��gM�c�m�i9:��ik5ױp܎�4��c��g��q˞N��<�؛sq�t��u��\���lp�4��K0�Yo
�J��m̕W��z-!��X�
�1��nZ�m��v=��W<�oڃ���݌s�ڗv��C*ƋB@&��jR�ֳA�ZX��<p�͟<R�t��og9��3]x�!�e����C�<��՟jv�Gg���n��sb���i��v5E���xT%-p$��]�+˨[�r&t��`CN�:��#�s�!���cٰ��M/V��P&��]�h�\��<���{N`�h�h��q������[�ղ�Ll�O<q��[���Q͆�J�]͔������	t�l�D���y8]ۋZ��xk���uc%҃�F�Z��ɍjw�����=uf6I9�4[�MȝA�n65���"����Q�A\� ]m�X��v��ΌvI��f����\Įɥ�
\��U,qr)0��I�1����h8���e73��fw� �������-]�]'�g�Nݠ#n�s��Pe�6�p���L��svt`Хq1i�J�#�.��ɐ����<1�F(�Li�F�bI2{ۙ��]yn�+\ݖ���V*���W!e{/n�qh���zR�j؆D�A�e��{�ny��b�a��94�a�$b=�)j�ز�pؠ܎���l�����^�!y�׮uk����e�q��Յ������s\˃��G�|����{y�q�k�����uq�:���6�v��j����ݺ��`�ǰr��[�f�s�!5ם5���mҦ��\��rl����>z��n����n�5�y悷׫���1� I�y� /���<X=1���s�N���/����rq�+y鵽���La���ab�La���9n��nM5yۛj�zi�԰�b�h5ѷ���A�s;%�X9{zS�\��N�Z�r˕l^�wwn:�GYZ�%Q����27*ֶ8���@�u�Wf�X&ar���MՅ�$u+��]6U@�4c���	��8��\]ãy�nÖ4�;9qm�c�"�b������r��$����0�n4�ƺd����
�ŗrn��s���2P.ȍ�e�m��*������4N)D�&0F�������]�������ۛ\]�:�m5�]xݫ��Q:��㹶�a�A]�=��k[75Ӽ����������\�t^:�n��[=�������*6:���rh �a`�hP�Ku�v�.ݷ/�_Y9c�#���2�vA�Q77h��6����4��y9nU���t�8���.-�Ǘ��78�X-�G6iH��Kf�����BF�-u�:��a�\.����lCjC���>6;�4�A�]�Vє��p�xfۜ����s�u\/t�^.���ڤ�uurgF�#��]�Y�ts��GU�nn�	�+�W���_<����8�r�c��9��Z-�QS&�a3u��<Vmr��3R�#��p��XH�bJ�k��f�60��\�esř�y\�v×U���0f#,]�eV�uɞ���YV�Fɭ/�\{rI�b��j��^2�ֶ����#�'������sڷk���Qv�Adȥ�x����q��ޞ�pD�5Z=v\Z8�s�ַQ�P���3�x��\���m��v��}�k�U�7!��nl�:��f��L��J�8��b]m�J���"[��bҸ�H�v�iD�&�֞5��}n�+Z67�4��5rַQs��֡=��⋛W��rV��4��qShǁ]Ů�J�lKrm��9���玱�]�طhj6̈gJ٭j2�Is�]�61����4У��$��eLf���l�΍�zU����6�e���ku=c�VL��_:�}���a{�;�o�$ޓ���:�ŷ�6�5�θ�C+X��n]um%�*R͍ڤ�&��Ǜqp\��+<t��Ҏ+��P���E���%����%�Q�ُ��3�ѥwTN�݇}�S��P���4�9X�����[W1�y˽א�2��u�][�{\=����vW���X��<z����ؒ�x�[�qu�l�B�%�.F31tu�5�����n�ղ�H�CL�aM�4�o%�v��i�6wF�dn��1Wl\;�wg�[�$f�`ȸ3����)]]���[Z�m�a�||x��^W���0�g�u�ʯX{�۝nf��Fd��f3"]��&m�M�Kh�UG[�l���R�F�Zb�J�GH�n.v�xׁ�ٹy���}�Ɖ�-�"<�F+iK	�
:��b3K�ɥ��#n¡v��6����+��J]-���7���ܔ�t�J�y8���/�뜏i�"�Q��
��c�ڨ�6�d�.�f�s\��	h�1�b��K��L�sL)�h�f�c�)����p�,f�Y�Ԧ$�y8�l�,���N��s,p��<qZ��ͮFRtN�t��4��Z�\�22�5e�0j-���T��޺�]f���f�x;v�����/l#O���Y��c��5�54��A�]5M�[50��F��V��B��\�]=����ڲٮ�B�`洕�@��v��nؖ���Qօ۳l�t�F�ك�����Y^�vDի��<�t<�q���̈́�%�*��#��7E,%��k
�\-IfPь�1�S����&cn$�[n�;燾������gh5��e�f]c%�kl���<5q�I�n#q��<]�mW����=�a8�,d�������u`�5���;L Uf	nԌi��e�K�s�LEF�ی�qƻs�_TН^�����^=`���K%׮��q��'g�����\/[�f�m�Ҭ�x��v��Z=z�=g����:5������ׇWn�]}O?6.�n�mlr���٠k����sX����G��2���0��r�
f��E�u��ڸ;EC��+'#4Ķݭ�lvvS6�9Uv�z�FM��s�(j##�v$���C�sZ�;�6���R�h攵c6q��y^���\�3�7f(qa0Ҕ].V�4����"�ps��F�t�=	�ȅ�GAV�{��a63��V��e�F�B�Eb�v+�a[Puy�̰��=g\�a9-��Llڀ�[b1u���[	�X��U~���?������� b?��i�E�E`���5�#7Tŝu�7��l�v��%��������f����3=��	y>�1�D�xB߲�K�+�xS���ȕ�ӽ�"��kf!Ek`L��Hl6.bb]��YsOlB!���E�n&6m��b��hdn�$��5���UOô��R��~^�h<�-���j%<�ڐeb�H����aփD��5��ǦSͽp�\�u�A_tM����Rȏ�$�M�j�F�v�o�q��>fϦ���^�{}?;�E��ْ��6�*v�Ӑ��pb�L�k�E1��������ۉ ���d&/b�9�}��Ǥ�ΗLs��3��0D^$vscS��V-�C5�U�"}��ÃnTY7n�WG�-�གྷ��]�9&�cӵ�:�1J�6��<�BnS�n1�Ek9���.�'ٽ�d�S)Q��k��1����Q^m�Li�L�i{N$��`돦�4��O/L�w(�������$�"��$�Re��ư���}�����B>�K܆7�/zj^��^qs�.����ogݐ���)�MХ�2����8�M�_j�h��= �o���8�8x Gm�,{�n�uY2���>��I"Aa-q�%�
$�K �=f�[�����>��"0���еq�!�G,Ld@v�;'�]�L
n����AF�g�q�Ý+{�{�aXg����3.����rr���T�Nd��T�F�Q���6a�.�����ֲ����V`�-�A�YGvR�N�Qr.L��2y=B����G}��v�[�4��Nh(��'ݓ�ݝ��X����{�wr��w��\U`�e�0�j��.�7ZsZ��(��}�TG��t�M����n.�j�юq2�G�ƛ��ٝ;dEm;�-lT#W/ ���E�1y�Ʌ!�8�F�[}���K�����%�ٽnh����i���bE��$J9!$e��^X���N�\���]��g�q��9�pjǛ���sٜ�P������d&�/�U`��Z������arWxAw7���Zz�X��.�{�gr��Ww���w��o�o�k��q8E�a�����h�_�/�����M�-�*~$�uХ�w����{�7��ZgF��;�٥�e����Nz���,��\x;PP=��*uy7� =냷pbӔ���x���̙�2p��]���b�X�O1v~��ܑ�r���B.�o_!��M��ʸ�4"18�x�B��ƺ�P�܋z��s� �(����_�B�*�/��^�7a؉����+͵pW�ヱ7������w�ꮃJ]7�� N���H>��@rs+)\�
<�K�vZi��r��(�$M�ӧ�/�//Lk��K2�gk�sI��ۋ=�s�}�@��^�}s���#^ �g�[�=܄OJIg�ǣӹI�&�K�tوn���>;wr�۔p�S��"�Ek�����x1��3X�{4��N�$8��Qn�e��Đ���W��8*��o��ag�T9b�@+��S��w�6��ؙ�.�K6����`���
Ay��݂�Y6�A��r����roxs[=���F����;2�Un��}��F�ݍ��I˱"H���αA�0ݚ/�/m�b�
ȓJ��L\,k55��A�\�[���YqR$=I�C��jfͬ��Z�Z�TbTƷ8 �/&�Ӭ�PX.6��G��|��'h�h�3�nN��{@�DΚ��W�:�&IY�{ľ���wf.e�~�	���`A���QU������j�(�R�$�cA;�p�O,�%�+��(�=�R�o��%��i숖�V��B��������V@��/���x�b[���(��8>Ú������|����v{+�z��*hbFհ�����Q��ÎЧU�0�(  �!�1Cu�)��y�0,;T�hZbt��$q���nf��E��YF��B�M#�,�g���R�n{,��y����Q�%�[9�a�����]@��f$�CD�Ysa=�wLƩ�l9z��$��b�c25c�W��,](F��F���&��۹�4��X�o��x��Z��3%�89NR���{��;	�C.�%I�Ǭx��g�n�����T�ٺ�~i�@��[���O&n���A��_�xNsnW�/Y״1����ŷ'\���˷{#zf]ν߷r5���.���_-~>4��l��M�e�/j��b7� ��xq�%j6�!`ѹ�B�KN�I�y?bi���~S�ȳ��˨���H��ڑ�qjmPn�r��[2�Y�5J�gO�{3e��Yq�
�؇�%���d�h�*DL�5� $�++�r~�#��$5��#�!�7RI��6sQ)F(+n�np=�7���Wb�_�.����v-�~�κC"��P�d=ۜGg��w|�����I99�h�&DF�q�H��!P��e�~��xy�h��ǜ[�u޳G\6'7^�B�n�7���R+d�����`IN��Μ�-0�FV��"6�y:�X�;m�<��g���orw t{;���u��8,�+1����������_�;�S�����#Z�`~�fIØ�ɮ����D��V�&p�f�d
�6štUˡ!Ċ�F��|F��r��ɐ\~��� `t�gH�o��8�<�i�`GOP[�P�jU�]�����AC�.kM���@�� ��>�*<�.��qgiǎQð`ʲ����٣��7U/r��ئOg~Sp{����/4Ǵjox��&��D��vv�ڀ�_�Ypnvpa���7)���k��9Ͻ|U�m��Y]�n�,�Wn�7��:^w�+vgQ���Ȕ)�UI�җ�g@�~"�7F'�/�r.��ȁ,I�\;���]��s���=i��u���5����a��p1�|uyJ���h(Xu�f2Aڨ��w��Ѡ�۩���Q3�+�����F��h�.�7�z\�&��#}�o�Jw>���h�}�q�=��<�)�y�Z{{�g{�7yՌ`)�+-�O_y�2-Yr���UnAOx��ۼϑ�����������O�,վx7�o��۹�q�2�_u��`�=�T�އ/�K�����hI{��w�aI�鰮�!�q��Oe ��/A�u�@�X����:��Z���R�ǵ^��a0�*VB;�e����6"t8��6�Ru��z\�{˹n`0�|3���z��r�Z.��Jt}�i�T��csپ�ܨ�	��w=�y�Ο���� �ҫbVU�,D���.�7�0�z�KQ{7��xK�2`��^�����.�o�ES�$�&�X�d�Ά-�QS&��w�ʴp��/hyP^�: �����b�b�%�dG��5���.r��P��x�<��7�h�ŻC�7Q<GQp 39�ه��˞��2�/`�[����.m8ِk�n�c��Z�
7f�h�5NBi׾;��ͦ���LgQvj���R�T�u���j�m�e���@�$7��ǃo�i[4����f�K�Y#'%�;)轅-��iX���������0�l*��>Ď�;��s�3Q�<��������	j�>>6�2�-��zs�y�����F��WH&�j�"e���x��8/f���A�7�č��?y������%B��
�Wh�#1�:&�EfhZ�l�.U��J�)��h��f����Ɍ�25���� ��̢���;P��m4ZYj�[�hŰ��D�hvji�E�C�J��^�4��zw������1�����H�lq�n���Ӈ��d^ka��6r�B�.�[Ksq�r�[�����S�����6���Ƹ�X�ػ^�nH���E�$�p�y�.҉[S39�����j�r��3 �3q�{�=�M��<��px:��wn�2�z�a��v���OzM��F!���ǻÞs�/F�AOz�̶�S�X�J��N��^W�P�{}ԣ�n������YKyF��,#t��Ef�RuV'*}CLB.��TPD�G�|$y�Nҽ으v_y1�3i*ڙU�(idFf��uc&��/r>�Z	3O6�TN�?l:
R�Sp�����P>QUR���mN�[�r>����q�U�Ř�~Z	:�Z�]�O�������ёu�ٻ�R�Ww:���3�� O$�}/~��xW���|4&�X�s���?�#9޽��ie�9��zT��	|�d{;o��ղ�g�r����i�b�P,��7Rup��X�b�ˣR�ᕰ{�.�!�@�������ōt��"Ј8�!�Ȓ�gB"�m�H��7{�>�Mu�Ўyi+x�{��@�nȍ��q,΂/v����I^��Q�m�L��d?� �#.���ӉIM�]��8�>�(t�M���+��`i�d�qK+�Y����<kb�
��h�3|�|�����0,�|����9�T@P�UeVD$�.rX nOK2!����
�zl�62F�1v�+q������������p� ��]me���(�dZo4��[M�3���xMݧ�z)���%=,�8ǳp��|}&tڧ�[����������ȍ�B�{�n��b�0]��U�d<�6(���d{�ݬ��eH�D&T.[�Uv�yU��*"r�0T,����ȧgrİh��o�4d^j�a��
����#��H��?'�w�kVWn?s�:'��K�ҽ�'_,!�(��hOտ��&~��0��]{����}w�f!3H��í�m�y.^do�����^�O�Z�M�9���
b�;ޖ�j>�Lygh���J2�Z����43po`�l�Ѝ^]�Zu��v���poj�|�}}޻��z�+��i�d�PJͶ��s�%�_���1J��Z���O��'�s��x��{`�L�<ȼQ��<�y��{�c{��w���m�ÕU�|_Q�#�������++�AE�%��9^�i�ê���Y��S{���v3Ӫ!<>�������Wg��w��X._����R3�)�״���hAQ0��7!���3��o��l��Z�	�xb(ycU�|0�gS�ZA1~��m˻�����"׬��3�pu�UTq��E���M���~�*z�ܤ���{=��W�3���o�) V�=����=��{�H�7pg�myO�y�<?n'c�s���O�� v��<�Y�=7 |MT����G�t���F=�Ó����׾/P�}�N��X�d�qɘX��z��ޝ,��h��+e�0۽�J�{����pK�1x�e<J)(��s9wy���E�7�9�&��-g��_�N�[�]�:'6�~�W���G��FbOŊ�xo_k���L}i^)�@�wz�e�$՘�)]�] �-%*�+`���8��$[U�y�B���2����ֲR�ů�\�3��yLe��F���{�~sw��Ew�U=I�;gʼ���vx�n�7���ͽU�4�1|�M��Nz�P��0=ѽ�x�ǿ�{)Sy�L˻�[��2+{y۽�ek{�O>"�����`�5'mT6������e��mn��y�~X��b㝨��_w��e��B����y]���{+c��v^&|5�4��Y�cs@A�)K�ҳZǾ��X]�ڗox0E �>��ޥf�':�����"�3iǗ�Fi$�E3]̦Mm�n�s%E�@!��ܟls�c��}<݅�-���|0;���9W���-�E{u&p���k��	�o"ݷt^�{-�`2-뵢��X�Z/n����au�\k`��!������7'�k*>W�[�u�yȠ[@Sw��n���y�|83�J�w����^�O�gN����:�s]G��\���byr����:���������-A6T[3h-ׇ/�z�Y�;��jl.(\I�J�Vr�|��9������8n��f�p�������TɻP�oi��TWz/[��Zi��љS�vظ1��#$��[�[ ��������ͳ>���s{u�����J	��w���[o�|��v	��F�Ad���(m���'����vhջJ����&���0�ɯwl���G����Pz�#��-T��M�f�ݽ�l��O�Q�>k��,�;�l�,�#�ҧ�˾ӸϽ����C���t�nE�R�Z�������l �l˰�2j���5GL�۽;�-/M-ɒZXN��#_�lz�bY c�</�n���^��qĈ�K�2���V�58A���I�͈�P�b���X�s�$KbZ506���  �s�v�wϡ͹�t^ɯ�9T�Ų�N�Θ"vܮ��>CZܞ�y��A�����=�������LYkiQ��Z����[y4�+f�)�u�u��7i��X���r]^V�K���g�m>Qq��V���-Ao��bbO?>3���4�Ro�h:x�n��k��H�x���ߋ*PH�W���orH�=��|B��c9�Ӳa\��)�un�Γ�j��l��ᤧ&'ƂMNP3pJ�sfwhܜ3˻Mlգ���x!٣r��mӻ/�PA�?h�  t�}�W�;_=9��H����N{M}��'��V�l�Ƙ��I3�{�9�Xnz0�q�tj���I+9A���KM��aԑEe�vv�l����~s@��8=��������:.]i�<�^��<���?vf�X-Vňװ/b\�L�Z�/THno
3��k�^�KDyD�T�@�UVRb)C406�a���)^0�wVK��%�G�9] �ΫK���p.���UKә�\�^;��v�fv�nY3k�y�&| �Y�|� !pa�\��v]U� Q� X�
Լ���튩�5�h��YN]�΅0�:u�٧"�!kov.����t�[��{-��՞�8�� 2����}[4�q�ԭ�;۽��|^�S���ާ��E��,�x���e�{عf�:���wi�Sb'	N첦��5~r��=��$ B��e�J����f�eH��]�{��t���{=�^I5�SnJ�P:3}IAFxQ��j*��
w�2�Jܾ�k֪�/UL^ץ��Y�5
�,����Дǂ�{x�Ѐ�ӧ�N�]���=ӄ޷"u�j.Ϊ3Z*	J��R�����]����@�"���
���\���g>��+#�tcBB�����WJ�a���M��t���QQ���b1e^~Q5�OK^w<�Cۻfq��O*�ķ�-[Rv��<='�ۥ�0�t. ��=���4\ɺt��0��˄=\��1�P��{@[������zΨN���m�;
���Yu386!0L�^j�R�]6�E��K���骫��!LьX�r�4
l�l�7MEiP^�=]k�Q�{��1�fj#��c�n�`ZF�e8�y�E�c�wD�ݝ��d��c%�nwpr��9�9��^�!�=����r�7R�w֣(�QyYv�����̈́bkT�F��FAթ����Ҡ�N���mj�L���š�浫���I�� vuՎ��J���}ϮJ�Ϟ�;�xcr��e��y���{�<��`[n�q��W�f�hդ��R]�d��Uٺ۱l�����NF�A.���a���jPlXטjՌ#�o[s�l�u�g��H��9^ܞ�|n/E���cl��n�NF�Y��!D.+��6e�n,t9��f1���X\�S4sG��Uגy�rVWE�9�Ւ{m���͖����W4q���r��Ȼq�G7������n0��^��H�%�V�rF��k�X�b��[:��i(���P!����h�b:�]��v�7O:��u;�Ŵn�F�hL.�+cL�Ȋ�ʃ,��c
�jCm4�iB�)�eH��qWU��P+s�KK���w-l�,
K]�8|���m�z΄�G�����=��r�ژw�lu�<A=6wg�oA7Tk�3m�n	�Eԍ��um�C\.�V�[�J�"�.���N�m��>:�3�ڲ�mr�c*�J<�SU6ƴ�M-��1%��6���[-auK�c�Ky�ҫ��f"�����ή��w��!t���y�M���cP��J�c��j�n7f��en�[R��t8Y��2�.�����	s��8a�Vm��yE�Y������sr�zf�p�E�2\n4��ն�"�+�{O`�5q�c�o7��j��WK
YG2�h�ks�i�N0�)X�J-����uX%9.�\�����N-���Q�7�?�,7|�GחLT�T#�ͽ}��;̉������4j�Fq�7�#'���D]촶,n��8M'�5]�Fј�n��C���!��~�}����D^WZ3�������><�#V��'��Q�b��q�E�s|�xf5��{�q��<���45k7{}�?Dv+��D�B�7}��y��ے��NE./�hZb�Ő��0�ot��}7L���޶��-����<w��_hC���!�-ƪ�q�;�j���}��.��<=IP����oo�k t�f�43x�:y�k7b-�Sl	[C�)C�,v��w�V��U޾���9Ek��X��SV�R�Șݸ�0D�lvW��۷6Ѯ�C�`FX`�z�ꎷ{鱆���sܱU�`t�<����P�݉�u��hl�m���|!fU��Ns���;���Ä�Fn]��� ��h��Q{��R":u��w�[��{�ؾ1Ϫ�D��1as]J钪����`Vp��9A\�Ѣ����U[&掠+�}ʸVK��p:�
No:Ib�rS���S5��tdMo��n.�=��%�5�v��z7���\�ʮ�Y=9�i�`]�80�}g��'@�GOs�q�`�gr��s��	kb��7[���4�s�X�v��-��j� W�tj�]x�̂��n�4m�v�)���7iUX �J�8g��r�{�{qy&zD�Ͼ�c�I6!�e�"�jS�_�y{���dk��{�^M�;��3{�,}�`r�;e��=��M�"�C�I�ް�$�<`]s.*�����n�:w��mb�t���yF��τv��6�����Wq�d1��br�V{����#���t_{���5H�ۥ�G�v���id��뭧,E�(٭inx��j�����b����*�9�ׄ�X��ݑ�dNI���OT��Jm1S%&m˂X6ch�V�E�:em�,�je��`KbEjq��ԍb-��uhX�s�ZݻG/W>x�n��d<t��B�\d/o�]:�`̫���[V֋+ڰ[0T)*=J�hDGedr�^ɭ@�!LE�
g.�����~�y��@�V�ʼu�����W�m+�r�g*��*py�7$e���ڙ��ݣ��{Զؑ��}-Ҽ�=��!�<-@�K/<�t��;�;��*�
h�:w��`�-��VZ'�D����)���,�O�V!�W-��C�&����Zܵ���$�suډ�����t M��P,��#u�:.Y��K�+"��Z�z�nJ�#tKuxEϻ{Tғ���^S�5B��d��N�
��5�꾑ӄ�r��:�RSnj�k�|��&�P�����Hb����g�^c���T����7說�,[����:jX��5T�Ң�1��s?\B�+T@�([���єk�Y�!�S�4F�v��nI9"8������ֹ�r뮠Ŵ�XSd���A�h��s*��M�]�~����X�m[ߢ8#���i�d
:����&:q1=��A�FM�f_S��i̔�6�nM3�8@NX���*1[�or�~��Ǵ��.�}���܈>��������@aL�Ɣ�_��Q�g�r�.hfIV�XS���cOZ=j�L���u�� vv��R4��^]N��R,�~�z?q�z���z$}�}�N�d��Щi�Q�uC� � Q�G��dE㓨#�Yʗ>�0,��U�5:�}�<�Q�;�QAU�%�LP�X�����:FfS�\��[
b$��ߥ�2������t��4�<�]6�j[n�Va;"�(_^on,dQ���x��`+;8�T|}�}�
�,QB��m\Y�b�5UTJԇ4��b����N�!/���SVF�سo���gk����&��w���o�h(6I�t�ގ�����d.m��n+%�6:��
��	>�����ݮ�S3|E�Q�0�M{:�F�{1ө[(ZX�F��]d�WPmP+)QL���KsK��|�r���\!%�w~q��(�o1^�3���	�y9�)�u��bY����!n�뵬�y��q:`���ҭ#�=H�U��#A���k��J ^,#̀����R|F�c�O^t��|�9�!|;�~?��t9�����N���_.վ�H�WM�o��/wN,���N��Ґ)*��GF/��&,Ӱ�|�l�z��}�sאf̴�x���G�#N��L�g��ܲ��e�KQ�(TR�TO�b�B��s��8&X���E��}���C
6#���I>�합�#�ֈjEK�v���/<;)������j�rb���m��;+��|q�Gr����'�p��;
H"�r2D��LJ��,x��J�ͮ���S]�qnn��wV�g{ߣ��|B�b��U7T�T��[��|�t��7F.��ǎޥ0�P �â�z��&/��T��j�H������ΐ���;�J��!&E��ݫ謋(������q^��xI��"�t�*|�JQI����}�֤-^Ӓ��f�E�)P�IWg���o/���(�)s��2�u˳s�u���Cϛ�'D�'U_lO��$d>sw�I�}
sq,젏	�"�x�>'��譠Z�3"�N��8��Tl��+�7�}�.	)��5Vk���s���z*���:SzЪB�d�$���ڳ�j�u��I�WZ�;�5^��J��_yj���R���K��޽�ذ����$i���ƛ<�s�rÞ&���:E�C���>�VD�+.���>���
��HŰ�=-�U5R!	��R[��r�ˈ���AV�A�"�����3��|~{���z���3���vQ#羽��蝟6�N�4�1	���z ���C�WWh�m�+"I�T驪�m��Ĩ̼����DX�w�qG\���r�$�ٍɅ�D�u
(]��ҵUO�s4��S1L�;�s$j^�TEn�fw�P�B�4evW���ZYg���pJϞc�r���lBu-����"b#����WadO۩���,��#�vJ���|�i+�],FnryM�@����ݳgJ8\��3���a�5>٭ha�A���ӊ�:}��x$_oH�,A�4m͡�O��ıIb��� Q�]B	 28Sf��~툛��>����n>��\0}�m�gd+!T��ܕ�kg<Z�u�yw-eS�n+��-��!��69�]3���H�*��f(Y��G��xɺ]S��NdjښǸ8��b(\Z���u�:ݵX�)�Ylt+13cT�e��w3cu=�:����|X�Iu�}2�r)\6�g����t��{cֻ\�v1�����M'��+���-����K��Ė���=�&4�;��*ﬡ6~]=�x���-X��������*�[� �X��Uf��M��T??�	���!]8u�$5���q�M@�,`�n��kl5�r��>x���{�n���p|Ē�����}�6�N�8~��Y�~H�"`���q��Y����)P	��33[�>���a
\=�-0Cw\��Y���D�/e]V�ԅ	|GHX`����R�	T9��:p_7�y���|q���!�foyW̐c��辰3�re���ۖ�ݦ�)�ޤ����	���z��e��>�ھ	t���l]��;)��_���,*�ciL�ĶQN���֖.}W����:��&$����i3gof��8A��381t���{��w\m5#f�fY���������]�,9�#��,�`s�bpQ�r�b���ʬ>�'��< 3�1h7o+L"�7>o� ��Of�M2#�����O5�j�U�1�I{��S�';�·Lu�I�@��ylNn�����z�	��C#ڲ�Z6"��O��F¹�x��Ϡ�Vt��I�ݩ�Y]x���ڼ�Q�.{����8@}0����W�K���6
��n�3B] ��;��M=���Q�؋���ћ.+O���qR��������X�0���B3E=k��Ns&,���1�
�Bi�GN�+5LI��3k�z��O�4�ÉR�d�3M�l)��!B�ߥ�K2���8p]}������Ht����iۘ�c]��jr�PS�MM6��+���Ǳ�@
���f��#�����|%X�E^�i���#��S�R��H��f�V[+mX�4�]Za�����[>E�{�(���s@�t�m�M��tV.���gJ�ymadQ��1�_T�K���eI5��Z@�I��컇�V�ZW;�S�'��:'��K�̘�K���7��a�0L�CK��	��k��<�SC�t4�a-�9,�s�ߪ�.��1 A��;�̒��g��Haɽ�(�z��@2`nEѹ"��j�Eb��������HxQR��xp�V
0|R� � �^��'!�B+�Ė�L�^;�g!��Nx��_ΏVT��վ�՝t��f���%�f��0.����d���Qdd�q^��q����$A�f	�˘t�r u}#��b#L.ް]����|�gDϱ��`��u3��w�.c����%˔�Ӫ�驄pɓx��xQ�38��HG�}9�d�q:@�T�����d>�w�����8ܸL��Yi��39,p�ԎV9{0;U��.�4Љ������:�nѭJ�gM�B�#���Ң	���2̟U���� ���	Y�g7�|�ȫ�eT*p�Tӗ�d�⧯*�l$+A�	��q�:p[�׃s�H���'�����9��>~S��F�^h֫�G��Rpb�^eZ�D�JS �	׫�%-j��븝"Κ"[�3W*Z*SuMR�݈�d.�^�ז��0�eO�Ѣ(޼b�����{�g��{<8�E	;#�I���(��;2r�t��U�������
�)×�`������>|f����\�-�m�%�ˋ�S%7����Ջ�{����<�n�r�u���"u�P]�	z�����Y5�� �#�KY�N���w2��T���2:nn,�����b�Y�)QD@E����|Ttp#-{L�.���jÓ�2�k��MW�tY�����Ջ��e�5���W�^�ZS�8}���`��B�J�jjF�Ӧ֖E��>��,�˝���$�{MW�/x
"�3���ǎ��D#�D�(�tgP��Y��I����΋]��ٳHgom�K"���/���b%p#�n̝:ڧ��T���0�s{���H�s?�=�����2���F[\���͐��h���3�< 4}�Hs�#�!!{]�L� +N�&Wg��)�ϵ��>ʚ�(�m�U4�2�����>��>�ц��B���B��3�D��%\i��7����Q�ىg�ȸ��:
oTh{;��1�v�zH�WK�7����������Х>G�D�=�g�	]=��i�}Ǿ���_���kߓv��.��#z
�R�KM���!Pt���Һ;+J)���ܴ&�UrF*�Ht�M���mgF�*'gE�s�u��C��z�zz�	4@5��y\$6�#A,�Q���6��B�[h,�x�͓hĭ�p�*�0*��
��u�<�n{n1�:�,�u�x�e�U�慄���]�,u�s���;v�=Q�i�-��9�G"���SM�c������2�c�W鱶N{;@9�n�uɭ�ʇ�[�4Ud� �	(W{J���
G����/����o�{t�UsdU����m�	n���m.c+����Is�7|���Ej���%��읜N��8gŊy���gHO���B]�
����Z�0������pS�.���H;j۹���>�Ȃ�}Ə����w�\�;��lD�B����_'V�.m�3��S�ϟv��Ӣa�k��k���xa�/:*P�4��!�r�*:.�� e�D��T��| C�����i��r{��iax�D�.(�eUlE%	��.����Ա8t����i����[�|G�6 �Ȏ׻af�̫�,�s�̫�p�z�>��j��ixbm���]IT۞�у���:�w��>Y{Ժ�<99��ZuD�V��� ��k�=LW�����#L�ٮ�_ =�i}M�2��F�gN�B�Qh�a@S��֥iiGys�xU����S�
.$��bMwnQG��<����>*��e+ Y�CO��33�M�]Ϻ� �L�)���$�O���a���p�:@����Fx[��j�$w-$}y"u��I��q-��"��r��8�'���ؑ�B�����p�w��B���F'H�ܱCH�@ZE��8r����q� I�$l��h���%���غH���U�%��q���	S"#���5�fG�k��L8%b�F`|0&��E'T���؅4D/�3zTQ�b��q\Q�,�S����ժ&Q<|χ��E?�u��Kr�)<=�������)�q��q�>�'�wz�i�0��˳,�:l��ݨ,�%���Xhe�4�X�&%��qnan���ܩ0�,��Z-���N4���f$G'\O	K��X1|A_w&����²�=JB�nWq�ݛ/eI}t��8�4�T��!���+è؁(�����)�:Y�V�]2Q�l;�g;�C��4�*��1��B*"b�$3&7��+�l�s����u7`Uˈ؈7nI���UN���(q;�_���{�ژ�����[^;:��s���}�z�Q3��}vv�D������͋h��y���%?p�p{@5j�#�\j�2n�1��;����߫�CE��s|&��M�c�D����|�l�BM���Y3j��7��3��*�M�"z^}��_d���=�X�/�x=���y>��ο,x1	�Kc��~L��<�@��D�J��ьW�y�k9�[#��Cy����ZZm�}g���cw���B�!�P��k���04�M;�`�����r�(�/O�c��֫{x�NGg��m|0]��?mƸ!ɴy9���Hc\$�q�H�����s^�=�����Q�EV�G�j��ݬY�4�/�z�PV��n���Hm�[�,�|�ߩS>KW�����=ǧ,�}7��(�G	��T�V��ɻ�]p��R�\�%1x����ܵV�Λ�]�q�+"����Z6�<�:ix�^�u��Z��������^+�ئ�Hr8Gq�˭{[�3qZv�e�K3��s�W�:m� �m�AQd�@�&h��oN���9j杞܇'�*e�Q(cY�jW�>�"p�xr��:��=s�����T��{�nU��}D�5�ק��3��tTq�	=������vl�It$��׵s�b��gc�����a���}�Ң�|O�|w>ą�U�0U��LQ�h��1`٪��S��2־�bch�{f��-Xz3p��N~}G�����t��y�k�����l�t'Ø�􉯲�4/��U]0��f/H�]032�1f��Z[���s�pj�-����L�U�F_=���K��?�m��m���~w�o���[aS[9�͝��b�1Q�DS������˛�ߥ:������ú���aEز��d��O)��~���Vse��b� r�����J�΋c�v�gw\��/Td��\"&���0�A�O��v�7����v�'�纸]��(�M��E�]�X��&9%^�c����Z7"����R�H�{�ج���O��t��`�'|
��7��lO̓xt�I���b�=�3xtUI�0�����n�FLh�p緓aN�f8�":9��U�
��}�������h��=�直ύ��r�̾�����HŶ4L�'�r���3�^�|�Ș֙W�T�EwD�o��t���1�^9��Vn�o�u��+3�^�=��f8z䙾���q�(Ԗ�S�b�ਃ56�KV��|������Z����Qox\���֕p+�xdx�:��e�љ�͗
�C��pʘ��Mim`F� �_st(�`�-E3LX�������9k��M�C��Ӊ[q쮫*k�vMC̽��&5]�#�Ы���μ��'�I�O�!�se��f�eC~��W��3�F�Jz�u:.��]�s���E�9��q�z{P%C��n�і@�Z ���<�;!Ĉ��c�Nʰ\�S�*��#XT J��̵����Sq�m��]wM�s�1�_�7eO��¨r<��9�J���6:���^�b��&�so˜��ܒ؜̵��ng,X��s��:�ᝧ��۽
B�qy)�ͺ�ȍ:��UM8���;ь��7:�q���*�j��ѣ#���[܊�&9��Xui���p�z�ٝ鳫���0��n��ϱټ�F�����:�Q�"-�:NSs�L�~�\���YǤ�~�`�mP�ϵ�!�����R�������P{�R�$L���|{m)B����0R�J�r^���m��)H�Hd����䧻׾��qƂ�fC}����������|{�����?8�6Jw�&����~��2R�/��f	@4��}�m7{9	�bd��I@�w��o0/��P'�dg�'R𯳐����kh�u����N@72�yܬA�R��&��Q�[&H;��$,�J9��O8���J����-`�CĜ�<�i~�Ͼ6�
w�%�rJJ_.�B}��u���(x�2^� ]�	]^��=6)̔����O3)x=����q�e�?���9���]A�t��H�%��u,�i��wfjv㋛n����w��ƍƵ��w�n�7����(�T�(h ��~��{��JP��dS����=��(C����;���1F�<�޶?	��)2]�)�b%@d��>�!K�s�� �s@{�����5���3�͉o{ٷ��=�^���2D��r�~{obR��)���@)<�!M�Ju��F�������$���@��	@�6���m7(y�j��$��!�CK�8���́�`������;�&C��������~��<ci���m�}��:�rJJ_a��b>��\�=�2]�H�f%�nDԝ���m)�2Cqΰz�M�hJ��d�����u ��%<%%*s9��]��P�)�2^�E�2�͸ݙ���CJ�H����\A���f��\	G�#��J�߹�M�}9
QF�P�pR��>����	B��I��#��{�q�)=��)B��rY@��u޺���y�<9�1�����n���u]Y�qG�r��>�J����|=����g.�*:DR[�]]�"��Ԍ7q2�b��ܢBӋ�34��ě�uy{��M]U���bj�
�Q́���
Z;�{�u(u�d	��'�����G����ߎ�S�V��}��;ﶔ�N@��R�(y� N���M��{�!GPqK���J�������C�%Odr�~��`�r�wߙ�'��@��P��&��s��n5�6��3sI2�e^��>�%TT�ۻ]aY�+�f�Ik�^��ߊ�\oy��x���>�-4�dS�����bQ�	����	�`��\!�S�2s�'��ѹ$�޹�Ɵ��~���;�
R�/Rd�y��y�=���"��(P��o+ji�40i�rSW��[R�i7K�Grk)��9�[C�� �+�
���)�`��'�}���/Ӓ�s��Gr�Cſ>�8y�=���)<�!�!8�^�l�`2}�i1$�$D��d�B���y��;���[�7��̞ɐ���(Q�H�s���Ծ���9�[�L��\���{���
���K��p�%/P9	�_woh�%&������)�_y��NHJ ��'���%%���Xf�Z��3`goy��_g!M�	Gq�|�d ��g>}�m���
����r�{��mJ����!7��G~s�n�2^e2S��.;���S�
r$����)~��9�R�)8�%�}��Z/�՜q���l޸�m�S��J9�����"�=�}�5���.�u'0䁹�M�&y��� kw�^d
]NH�)J4��ߵ�n�rSy�����/��p�ԡ�x�ҥ'�d)�)��-���k����:�����q5>$Q�Q����(�z��Ǡ �.U��'\z9� �,DĞp��Q��}� ;�r��K�ЈH_��ըvŵP�o`t���8Ln�A!�`q�]�.*V�ڱ���,ۛ]�sc(��hE�����aaf`�ԅiR�u�s]�1�T5��Ԍ�B�;)ݏ7�e���퍇<�y��������R�Ǌ�PѓG�=;i�N���۵�;Wn<��ږ]a�X!�%�X��m�+�N˼�z��DG.��Nr�EE�1�9���n��jX�1�
O�eG���0_�_. �����U�f��ې� u���y���/�n�>#��uʝ�^�C{4͗c�c��+%�-f�E����������s�����;}_w�9�2J_$rSy�}�����O`2��
S��(��|�[�6����9�HҔ���y�^�y���u�p	��Jud-%% u9	�����5+�����|�"B\���I�mp����IZ�́̔�.��:��b%)By��i�g/�FG�J�)JjC!�
]�Ͼͼ�@{	�4�I��������ud{�Ҵ��9�QǾ����L��0�Jnr
]fQ�C��D�
�ƨ�R��ݻ.Dx�(��)�p��_y���s(�%hh|��J����fԤJN$���0����b�{�����`s"RP��#�b�	C�y�� ����G��(��i(l�VAHK�RA�j$#Ò���%q���|�h���)�r�_w�l:��bJW��M�
S�w���7/�j��C��(�@�|�~��P�d�9��㏝�er�rj߻��o0��P�I��pww�<��;�����=�t�_w��\k{R�)7&Hw)���P%��=��2P.�!O3��'Ԏŧ�ν�����ry��.Gp%K���a�<@���%"Ry&@NB{���l� 2����Gy�Q�n�ٳ5�F<F[�3��v\[��n�i�E���9��b]��[z?>�}���m�+�'绾�������N�u9)�`���[��J��]f	@�w<é(8�}�׶ޤs��8�5FE%�9	�}������d-������}��<�����kj�%%(jr��aB�$-�ؕeC��Sp��r��}0�:�7���#�pCRRP<��ñB�f=	o=ϫ��n���˯V����,N�<� ^ۉ/�Y��a�1�S
 F�{�|(�]$y�F�@�pf5�O���>���P%�9�P]P�<of�Jݠ^�UIU�ۙ���M���ʻ�u��� NI�]��7T#��1� P���5�/��R�}�$�|��)(_ �Ns)�|����W�#��z��O3(�<�RgZ߹�(' 9���� �C��)�2O!�:�ϸ�Z��M7L�p�[v\pP�f �$���C%�rT�ϻ����d�� '%7��G]��Y��h����A����(ҝϺ�(�3�>͏����Q������^{�m�@�1=� ZOd���Ox�:��lLNO����o���������q���5 R�fQ�}���\����b�s�k��ٱ��%7�<@)I��/[��m�Τu�Sԡ�P���{����x��C�ę/���V�@��߇�t�Gs�M���$���8���0R��|�u��_g!u��;���47g�����|����N��Oa�z��N=���[�����;��:�R�x߾�Na���)�`%�d��~�����C�X�iB	���^�["#���ط^Nͺ垧��{�����:��W\:�޵�����a@R'2d�y���a=�������rD��z���
P�L�;���b{�f����u9%/P�{�(P�����m�r�:�9���IIF��ʡ��)�N��v\s)�b%)I���O����5�(���!IA퐆NII�b�s���S�2h59 {�%��&����J@�rSy�p�JP;� ;��z6� {�%a�KBw�(i� )�~��|g�W�ͯ��jR���%�>�Pu��G�{�\ld�iw9J�������\&�;���0~S���z�#��,E�1Q�*�ԩ�vmؙ��,�����_Ʌ��a�k�)ڍ4=� ��na���y�G��G����U �6��0$F��·��m�P��g"m��*�V`Uy���.����wz�9�y�m���|u���,W��2��2JV�޻�8w'p�%'��I�R=Ρ8�\�fÈ\�`2F���rW���p����	t77v��K�A�d��'��:� �{�hђ���fҗ��3�i9��%�{�S��(�@�))z��h<�޵��Д���{���ϐ�h���>��m^d��y��%ڔ��JE!��5q.I:wSwy�ܼ�J�1�\�%rJJ@޼߹��Os�)O$�ԝΧ�0|ҙ������A�qI@NBs��s���q�5/9	{`@d��>lؔ��B��)7&K�>��مFZ����8ۚXe2�5�]�WZ�����zm�97�;�����,E�������߃������ߓ�d�K��!�o�8�͉F��$���Ns�#�y��6�%�d�������)<׾���y��/���f Q�BRR����w}�%I��J�Jq��MRr��JT��t��Z�D���R������7��}�|�7�P�%�r��0J8� JN{�{6��Ӑ��+BRs#���?zm�P�0Jz�28��5s:���{��-	N�K�^dԾNJ��ʄ����t�Bi�m*���IpPI@�J{��@q)�5����/s���P�@d4�Bd�k�=���`����N�65�ɩ{��P�o�OP%K�����������{��b�RB���R*�i�&�q��nD|9+��(>C�)7&@����m���
:��Z^�!x�^|fĥ)5&C�4�'9��{����̥%/�	�b#��\���O������r�i`�}�ڍ�D9T.�|*T3vMԶ�'nr}�a��(���GM]���S{:KW5���mM�eMC��ԉ��j��E��ȱU��dRQ��ﴰ�߈������)˱����a�`W�*�y��>h!#�JE!q��p�"�}��$x�)GRs�)�d����, �)aԑ^���9��$ra2��C��~�%��4/s��f'�Һ�9�m`~�%�r@�0J9��7��}m)_`ʐ�b�	Hs&K����6�u+�Jp%%��'�΋���ke+�1���#�:����rD��n���ˢ5�9���M��;���`�\-������y���MK�y&�:� ��n:����9����:�J�0J ���=ͦ����M�Gp%+K�wﹷ�>LC�0J@��L��r�7��g0G�IK���`�Z���}$�ʖ�EZ���K�,"�P��By��G��մ��r��4��G�`�)I���|�����`�u�RR���}�z�[���S%�r^�9�	G|yϼld�����q����	�b%	�����th(���}owǽ�<���`�wBjJJߟo8w	�c�.BR�&K��-��Ϛ�"U�II]�����=���3�C#�9��-�/	�b5��IϜ������u(s�%CԚ�/~��?��� ������{�w����wy;��Qs��<pOPS����)���5+��M�+G]��Z��IK���#�J�$��=ͦ�{�!7���d{�&��h�SA������!�`�I���B)z��S��Rn��I]��Z�H�$��^��M�Q������S��f	F�޾IC��9޾�6�)��'�B�%'7��^u�ت��/L�=��vD_� ��=j��<!^C���@�Z>��w�ّG�ng�Ͼ�"0>�F��b���빮�²0�(kҳ�e��Jf<���>��fԖ���M4�EV�HJT[W'Bq���[ó�wQ���ɫ2�35�۶t�/!&�	���կ�wGL���l]��rÆ8W&�E�+�Vͦy�ZM4R���[����05�]�l�������e�ۊ���\q\E/l	�ShU�[`Ѷ�(�e��Y�:��2E�F3&��6��Zں��ǢR	���{�<�w;6뿅U�qQ>zP;R3�'`PӬ�Ž��z�T,ص����L,�܊�W���{�)֒˂�>%n
f��ݨ3Y��uۄ����i8�.h�tv��{�=��OµM�J���w<��U�$!,׵xr�0�*`}ݗq�ʃ�B�3y5�(< Q�$H��1���{��K~Q�H���
T$�HR,U^�`Z	���v���%]!!ɢ�VLsޟ��(y�1�Y�}�X�F���o����5J�IL_��%r�9MW�n�>��O��=��kx�]�������4yB4���EJ��5��e\/L��_����eJ�Lv��F>N�U0LjiL�'.�(���CKE,H�)����"L-�0nz��-�"�����{<̥��_.�9�:�Z�:�c�ʝOӵ�Sr�Ljқ���C�)#
�#��^��I X}�r�~��x/R}�����&P�5�de��Zgr��I�{���!,0�3Å���Hm[��+KtQ5��̹qi�����v)w�I�T�Zw�X[T���:wO��].҉�8�=<��%��I��p�bb;<(��~�"0��:2}��
�����B�6i���M��4���6��}�Sg���T����O��b?�-�i
QU�q�Sq�p�^���a ��4�I���l�*#�Y��<�>�.rC�vG%(�խ'���ս/#)����n�T���Ħ�!R-ړh����Ϯ�:R"(Y�TX@#� Y@Z�Ƶ�MX"�� ��)�5Q�2���.�W<�aCH�Rs��=��4�*�*��H����¼vk﫰� ��N��E�� P8O&�߅`!����]n{���B��I\�麧[�$L�9�UH��G�����A{噳!��^�c{�O �œ
+��䪃BB�Q����H�
�J���Jj[d�&���B���3�
���92@�<�	�8��ݪV2ad�P�wy�!\�8J@�ǛO�9��>ny���C�۾[�捣mh�s�nw�u��`�^V�pv�Ŧ����G�
�!@�UJ���&Pk.�H����a�Ļ���+˄l/.��� ��{?��Y�A{�$d��|�*AJ!%^	L�
���*.<�V*���LGb���i���%���_�WƂ��]�s�x�� �^�)�}):
]j_нo��ܟ�9�Q�<���b��o�j��g�sq[ˠ�o�z�Y]y�c�*�ޘ�.#�c��9�f�>ƼL�ڪ+���׽�$Is��x	�=n�()�sb���8���=��<���>ޭ�f�-�On��(���0�#�5���|c1e5}�8���i��B��SE�+a_��(���W��0�]�ES�ULV��W�!rW|��
��o}8 |�����
���� vz���G��\�V�f�u�٥�Ъ�v�v=TԺ��n�R)�i���R��Vr�P�5Y���u�55�lj��آ�-+���}c�@W�}�=��>t�q�eI�S�U�����*Ń ��5��Y�oQ��וa�'}���TW��Ӣ�H�^w�+������%xr��� E������C� a Ϡ5�ld��7�I՛秓ٵr�h��=u��b>��������GS�1R��������ߐ��S`�  ��"b�����K9�9�>�ƂM�~�룶*�m�P��^6W�{��8W�W���E��
.�g7�M�<���v����Ԡ����*d�(%n���!}�����GЏ�T.�v�}Ƀ&�=~�⍈p.|�u:�l���n>W�j�v������)$׬ۺ{J�S�/���ޝ��1=�G!~��쭥)&`��>���|���%���r_�z��F�W9�O��$-�UȷL%D��}��e����o)�C�t�U��]�<�sUi0��t����]�$�qy��m�Z�!z���_��S􂟧vy:���tI-r6��\�f\Nn��k�Y+&B�!5�{�N�Y�)=�w�)2��#�x�+؅}�*|PT�P`����P8�kpW4�S(��Z.+u��#�����k����*��D"c�EMg�=��+뮠8ݠ��>�`r /R7}�� p\��	��^�s���S�g����
�橷��r�J`}y��lߔLBb�8MA�`�C�-�=���f�)_��Us��� CHr��/䙳�;�*���1��5F�Ä F��0(+Uy��_����@�&����}d(}ت�ŕJP��R�0&�"�T<�(!'R7�ϯ�O��%uȀ���+ڬ��������Lԅ폇�"N3����k�1��ug��}���pYu'<fj��1�^�|����4>�����{�|^�(ӽt���zJ�Y{���B0l��!�]�d�.6�^&Nw�Ũ�K����v8 ��p�+��x�N޼;�墿c�~Yp����N�ώ?�;�¨���Nq���Sw�e�c��3k �*qC��r�ws��	\jI e�����?�����!�ߨ����;�)��0�V	�w��tk��펒���S���ow}�xok/�샚{��-9Pn���.ޅ�3�Q���^v�x���������H���I�MrC�~g]���!|c�K�|3�;�^:2�j.DX�82�e�lD���U]+�SP�U�X�-�eL]�n��d<"`�ln�Ɲ��r��;p�����e���َ�q�}$ow+�^ow�2�f[���&�n���8:3/n�)��?T��}
�D��t�9�Gmj�c;�F'f�f\q�#g�����dU�y=�����J'�ȳ|�5"f�s���-��i��':�{=~�>�%�LG���c�o:�*u�)P�6�in�{�[�9�/P�V}{�
O�z�,��V��ţ��tT�c��L�T�0���
M1�i�{1�
ʭ�	B��
�t��޸NO�G����G����k�ޥr�U�W��m�x�Q���i��Jct�DI�]WX�E7K�F�Q0g���3nd��Ov�}��3ٲ�X���:nZJM��_��J��Uס�<�)s�-\<����U�)�=�]�b��#�ȴ���j���_��89{��	
}�����q�����c�|j�u�u���c2(b�W�
�rD�&�^Y%#��*�h�z��T����Q�fv��cm����%ӻ��L��
"��2�Ru}����&rw��}��J`�w4�֑���6Z@w��ﾔ2߼�@�����ŧ={�����X-����v�o�^���"�3��{i]�H��{9��;�;uwLwkW#u1�˔��DD!0�z5�-c7�qh�=Q�i�`��gk\�Kc�]%,b�+�un�f�P����ʕY�4��T�� iai܆�c2���֭r��x��t'K٬��<-Ő�L�`E�ۙ�\����n\���f��9�+R�%���HhM��JhK���6b�.��B\R�U��n�\�9/5sø��ֻOgqͷ�ֺ|#;hS���tø�j�Iբ�}�ޙ~�\�ɍ��N=�p�vn=��s��nڎ�����}צ�t�z{n�@)9u7;>!yk�ؼ���lw=>�;����4Q�6a�uV�ڐ,��ٛQ�:�{��%����9q�ہ��ź�Q��헌7��)eRP�۬]H�k����eB���Y��R�D:��KͶ.2�E.p]�c��ϡhJ�=�cvl��Y��s���[�F�ù��+b�Yˋ��"k��upث�˻F�z��1�۟��콷��V$�-h��8���7-<��5p.��u͔es�Hs V�&��h7U�o��/|�Xx�kvݫ��G��g����Q��/B����S�kc^o�d�u�2�S�g#n��j��{"��3�8t=c=St����C馚I�n�ѷ��*��S�,�2�-5JSUڲ�<V��b��%qo<GGn:�K�tc�;���w2n�	)z�xn����S�yM�خ5�r���@;�j�|t������N�&��f�����Y��*h�6�(��׶��#lWm���Uth�Wۖ��Mn4�lk� �^�Zf�tf$T��xFna����:a�8S��ﶛ�"���Az�jS�;g�bzs��ּ�I�J|Yx2�b�a]���X8궹�z�n�88�n^����u���뙇l�F�Ƭm7`��볞l�cv㭞:��O�Cq�m�-����la�vہ�,sk�
��ƽ�<#�^�n�!M�N�7�����ΈB`�3(��=�_B�8Aġ͈����u�t��7(蝜O�n�6���D��He�P��ݥ�n���*:*e��/ThS�16j��*�g��C�>�٬���d~�U��UR��Pr�Ѷ&�Ua� Ƈ&��=J�&�+ّ ����M�\ �=Do{y�
�3�v��Wn��^�`;����V��|�p1Z0tE-�QJ�\e[Tc��ev
�-[R��e��9�b��gLݰDM�3�z�wqqMɮ���Ev���3�Y���T_�\�݆�0��)Nֳ�s�^2�D����6b:�!&�B3)m,�Z8�S�m�]������<h9�Di�`ʾ��l���[=rc|�o��5���P�����哬R�@�F&����|r���7s���tmN���V
���;A��To�c���C��l㌿B��uBC�ڸ���#�}9���\���jrU�����y�Z�=�vƛuU`���\A�7��[5f���vI�]qqn��[����n�'�;���h5���ٟξ��D�F�l���ʢ3aҍ[����)�mw�)�׀��I�C����	0�~vl_G���q|4c���� �B2�y��WdZĹ^R�S��D�oD�΋�F��=��7���aw�������-�j5G)�ET���J����t��#�j��аwP��:a/M�K:+`��S�b22m)Y�w]�7�"W2'K��0�Uӳj�X�Haĥ������wC���_b�R��1��YSm6u�ח�r��Z�r���ۛ�X�Gg�T�k]�t����۰yJ�����IA����Om3��pE�v榚��\�Yu�jU��,���5b7gA=���|�s�⭮���[s��}u�qhH�����1�S��Z����>qݻ5ݹ�5�����v5�c9�j	��4����Ŷ��A.C32IC����v�}��'ٌ����m�J�{c��0���b��l�����Ʃ���&��̥+L~��w�*ܹ��{�I�c�չ�
±jX�B��ڎթ�X��R�ۜm����ضw���io{à@4I��.�#��J,��n�h�_+��1��f�F@5��i~>
�}Z*�V=�zq\�����gJu�T&�-՜�3�?H��e��R�IQt�?_�>�V�.<�K�ER`��Y��,�j�=	
: ����y�*��)�(�˺s|+>E����q#�
�+u�]�O�0����o�v���)4�ɯ_qP!�Кw�DI��' ���6!`P/��$���r�JE�R��y_#�����d#姾G��dA=y��\�H�ɏ]U:	�N��m�}9���]]�)�=��C�@�}��$P���_�`�Y>PQ�S���A������Y�`�G:[u"��n`��lHVÀU�y�p���2k��s�Nj�{�}����uβ\���RY)m�Ռ���wyW�NJ�en��!*9�H�a"�{�|��4�&X*�ʨ�7S5ɛ��N���#ʺ_��30YA_��@�$V�O��������u>u�g�DsT_Y�g2a|DpV%b��{3}�j�7j{��E�|�^����}vP^�M�	�+�;%��K�����ͪ��^��1���)�
M�nn��>����#/�q�`�3����� ^8�| X'�e�Ý|�Ѩ�����׉�멗i�&{����r�v����OH�L����������Oݞ�+Й�gt_1�;e7V�6~>Md?{97$N������cc��0��fN�vEŘz�N����Jr�����蚖�B[�'�v�������^��CݘÇ��%I+D?�~w�h�±Ns�g�>���id��Ĝ�B=��M$�����&M��Ml��uQ��M�,Tլ�����m��(������-S	��]��gj'��yW���&�I�n�k��:)D�B����ƔA���e�����Y����%#�:��Wut���#��I{����B��u_�S<�K���N�wy_r=

(�|���}�뽥���u˚�b}9����a�v�����&�FI��}}�]d/J9'�����ٔ�^K�#�>İ�>���wT#H>Ɣ����a�������x��Y�0=��m<A�k�]�#�bnb���Lz�jfx	k�u:j���^�u�=`�n�m�,�&%�� ��n	V��xb)/>�#_���?�I������V�(X����%�ʩ2�t闢�D���'DC9��QF	�z��qGD�ec}(�:��(M(�.{�NץK���{:MIHU\����t����}��ʳa"������
צ���ﾫF������p���>�}2"�6�y��+�v���l����W+,�M,�J[3]B�G2˞�2ש,�f��J��t|<��@]���r����~��!w\���>K�����y��Tɂ�{�4�UN��T��7iܥg�9�^?(T�x]��R�J���J�N͔n^z��s8L	N�6�߀C��>"�%��JQċ��ب�_]I}��޾�j�|=�(�
NUׅ�L����뿶ddY���%Ԓ���i��5�g~�,�]o�V�g���>�|�X�Ewv_Ƒ������ФQL����E���f���K��8�xNA���`0P$v�H��餒��`H8Au�(xQ
�������N�o�χg{�Jn����-���i���ϻ=���#~(c�jt����5�=���8��ec���� ����!Yz����l�䮰fP��-�e����.眕yz֜���Jb:w<���	�j;3���X�ҕ�̼���:)�}���{{���f�L��X� �����Gg����n�˪Q+]�HkV�&M,+^J�R��]��ⅻ1��O�tg^U�[��+7�u�Q3LG��]x��O'4u���M����5"���m_� e�si�w��a]�0O��;�v�3�.�rΑs�ٽ0\�%�x��9�Rt�m���$��_zc&l�o���D�
{�8њ�֒2S���ޛ�3�+�}�V/ￏ�C:d.^�N���C��^���+L�����<櫞OH���Ţ�t\�$��(\�ÿo���&�³�>[�9t���e>���Ӝ��_f��z*!��0��ަ�0�Gsoj��(>ҟ�P��O������&W�D��_3��|$���*f$�!4.��E��fEZ��]�8�#�U!���Q,|����O���.6vm���F�K]�u�Yc��kp&�W]T�AŰ斳Pv�ƭ�,hR0i�g=�n�WP�9��Kô�gx���Gi+�t��q���kBE�]m{>\	֬JD�4�jugqz�!M�ė��q�/�^��h�-�4�;�/T�-��^�݌��J�ם����/�\�F�1�5M2�4��B����s��ai*�̸������j�n�W��^���{��Xu�8�ۭ�V�{ǋ>���28?q�p�A|_e���~R�l��=���@��Yi^c����Q(A�%]��&n���x�����ڛ�:X[T�V68q~s�NlN��k��	��Bn��O�ɞ�7��Րfś/��T(:פ�<�~ �d"�|t��>�7U�h�,�������n�R�TTяA��It�'lG��@8�7�a^0�y�(X/��5=����0��A$��x}'��ߥ�l%�5m�z�x��F�u�_�P4}f��5����@	�>7}��V{��[~�q�8%��O�J�H��2~t���s���Q���u��*��#��?}v�W/i�'k�ZB�ƫ�鄗Gw��b���/|��%T�*��w��|.�6Z����?(ʄ���|��J�G��oJHݼO��H�z!��Oڴ�ikJ�D�r)PǇp8�Kg{4L���4J�˝\n��㏮�����M����Gϧ�W��F	�Vq֋K��+y���T	%��Lp���Va<��ީ<�����m��y8B3v^����W
�Z��#�����9��(S��_rR��Ԫ꿱u�<B�TE�#ne{�~#�u[�x�������s�Ai���o��O�lu�h!_�zM��qH�o4A��Sk.V��+wMQ���FNg��9m�ϙ���ȰW;]>�ע�HQ���ʉ^T�"D)D��SD|{.=�����,�F;��p��%1��㦽���ܭ<t�S����wf39z�EQIÖ�^,򉄨���J�]�����Y���yu����O(��,7��;�S65�@������4ѩ룖�At�����? ;��)0!�}�W�)\�`���^���D��74�����H:
�7���Y�1��%�V��+��5m���rK���N��IN=Sv���YH���->��O>\@��1��W_xG�+S?}�޽�uύ�}��۽�5Ê䵶��>]�/wg	�?x����Λ�(�K���S�g�JMG6��_z!��,:o�*��D�h�E6���ȳ�����V$�Ϣ���ބ~���qɱPWd4��E@���^+H:`n�H����b�D���xH䀳$��`�U1��za
>E�4JY�)�fL�5����4R��$���ٛ���C.�\����ƳX�3����3r�	f���ىd�߀��/�WF* ��U�%i���*T��R��b|V����zJ!3�W�礚.���zY���u^�?DJT ]���aQBі痾֙.��$M��4��͕å�Mi󕢟%""(��߽�ץ3����.P�^fϖ���zU�E���|C���� F�[An���liRL�b�P�0����K�-m�Қ;~w!���j��#Ci2~.�Xc�Ί� �&u��\���;Y�M�MH̪�V���!ɞ��@�n��mլ�>c�w���C;�����?J������eضo����� �$�F����|"T��	m*�}aI��{�Pu�GKۚZX���I �A�{G��߫k��C9i��,Q��D%�PRz�*���L�<|�E$We��q�8���O��W�L/Qn�$q����M���'�6n3���b<�*� .��ے}��	���QC��>��.�VLT�>���q�_RA�P&p��+ݺB����A��0j��Jb2���聾����+�^�'��;�����Y�%�
Y����y8w\�P��}��*����n$}�o z��FaH��̘v�g���R��+�%BN��X+�Ǒ��}�w��>7/�/�V#н�S'�Jcx:lm�4r���n8-��bgl����O�����x�S�@�m�����e,�E5d��ۊ�����خ~�>\��9����凌��E�S�l���U�䐒�-S필�G.>Κ�BO���G5{�zϙl�^��|!�������,��l�(W�K�g�{u	�B�K��O���|~�K.��<b�
��V��HD���e��J���(S�����w�Q<wxW�q�Rp���ȯI��|<� Y�6}�f��YP6;�P�ȑ ���^O	-�,����"�%�믽W��*��,,0Y�Jg���? .��T߀�RI������@Yr�tT���5 ^d�o9�����8����o�z���ߛ���߫��sֈ%=x�7h+�Q����u`=����s����8w$Í���5��	R�QKu�8`7X,����WY��r7\�55u��y)yF�C��%�ή��@1`v�A�W�x������=�kn�t�[���%� �`�H%��q��TSZA�[�i�!�j��^9�OV�����N{����\/;��:�&x�(ԫ��Y{�4�ݠ�)�uq�4CN�P��j�V�Rq҉������-�
h~�y�g��6��OL�#>|��Mv����,��ɳP�Y�WQ�8��h�;.��L�!��z��Γ���9��!���t\�*�v^�,"��j�$D-����`�s�ZpR��?T�`4�LK��i�8G����O$�B\�5>����W�K���)��}ʸ�$�*"8h�3��U)N��uZX�A�0��t\;o�g������w��K���
�8�(ZO'/M>��n�U2�楶^���DD�fg=Mif����^����i�F(�da >Euen�ެ�}'�_��r6\(���a"��Ҏ�;>P�Hox��M�NPN�5m>����Ը�#�b�7�r�E��0\�sm»=�0�L�T�i��J�%�]
����]]�T\d�z�]n���,^����ذ���O���m�|���D��
w����%΋���7�*�
BQ(ʉ>�[(3���9S?xy��*8sbyN���^���8���)��₸�pq�24�#��}5� >��B8C��"H��!��v���pv�q��^b8d�L�������~�w���q�4[�)�~����{���(/I�3�@�sw��շ���G2�~�^���/����1���4LS����_�U
�G%z�'�;8�l�Z�&˺���|���ݳ������FM�)�`��}n=�iû��^�gӈ1m/��\�6��KFg�LG�a�{;V���7�5y<�|�x*0�)���M���\<H�|.��\�0LDHID���k��C��_�'��{�\��S"�>�>��Va�'���Γ(э� n�%
	��	>��p�h�V�K!cs�F�n��jc�X�աcT�۞���Xi_��`;D��s_��Ǆ�������a�Q���/������)��/�rU��'�'�|�>{7�&س#F��xN�������a,>+f����_Ef�\�/�QMY��u>�}�Y�d}��*�T�l��/�'�V{�W�,�,4b�(�~W�X3h꼢M����� ��!+���h�#{�d�k�ޣ+ )�*�%���4os,�/֥�Y��+�r�ͦUɇ�Ӎ�K9h�S�a���sq�=��쩂�6^��l�l�'{]������⹦/X�y�ocDO4�{���[��{���w�HgR�/m�w����+���q�:v��V%([���&U�W5M�����I�*k�>_k\�}	C~�g�'{B��#����r�(��軴�t���`>@���o���2�M�/T!�^�\O���f��s��/1��|������Ͼ'�̫�g����i�����׍r��z�6ɑ�F)��s��^.�"�U�m�R����E�T[�c�W��8��[l�?��Jo�iQ�����#ڳ���1��}�*�x�p���K9��QuѵNw�nj�Oh��;�ځ2*j-VΡSَwJ�n.��}U��u�1�p}����Ge)�'�oJ�k�)�]���.v[t�����5�0m���]�~���j/_t���'\�D�����q���A幻	��6n�����u�b?	YN�x�_3�`�F���v��G0�vw�m��٘��zos���)w�Ј늓ѥj��V�)�e꧆�J��IkU�lQ���^�������9ٮ��-@-����'�w[}�G.��@�]w�Lt�XF^������c,�ʜ�
�c8[��v](����ȸ������|J�xU��e����F��q�J�wP����#���Q%�����5��=]"�c��&��J������Ð�E��ˈb��k35�ˮª��hJ��9oLvEd��շ��3�#�R܆�����,+�����J�ƆNs2k_���Rl�ˤ��.�Ι�:�4��\��<��F�a�[�h�κ&���sa�[�I�K<e�îH�˨�ӡ�p9�f�}'j�vs�(�!n��5��FS�����o�ĳa\�I��p��^�v��ۼ52���r��d7��C� �q��f&�:��Uu3�ai��=���V/"�Of���[�c*�P�S�xX������og+ދ�G��˺��;5�s�XB0���,*�ڋ����j�9w`�׮n*��u��/�0�6��b�~��V��H�3S�י�m�f5>�����KbӘT]�XxtU�s�Lk�_H���;�W�_���#nP+�랇�Ld�A��9N(�R4s���J�+v{7w"�dPAaɥ��wk���8	zTDu��(ܚ�t���f�Iʗ:a�h��ֺ�:H໡K�t��Hv�(_F���tC�]�݋�N\���v�"��n����Z��6�6�t	��ڵ3ݑ:��nT�U����ɂ%�d��q��\>�%���NT��f
+`=�)���ӛ�q:��=V�8�L���rh�H16]y������a�~y��-��Ki��vB�����Q��T��˻���F=Rj�ka�����A�m���b՛��U\��!�@2�LN�[e���Lj�¥�,Ӌ1ɗ��c�r�ήg�A�zE�����W�P�/)�n��Z*͉��Gf���0�^S�vhED�w���W�7�&���y-������[z۫*-�U���R�3bR���$�nX&�T*P��d\�jJX[4����s���Q�HI�%N]���I�
R�&�fUꜚu4�C��Ksq�8i��PH����^(]�����;�K0��v��X-4�b�~��EF�p���)N�3$�)��ŝ�����G�O��,�ߺR�z���/��*֗��O��V��9ZG�I^�*��9D�UU5CUIe�e��\9�Ff�%SY`n��5Ѫ׹�)�b�JDH0���\D��0��g2`Y�8_U��r�Κ1K�����=��+��Ĵ���S����Ck��*�]��Z��8.�o�p}^N#�]4V}S��07�'�D�)��\Ejg3c��Q~>�'ܰ���\�&��/
Jᵟ8��7�����"raGO&ib�g�w��Mdʪh�,9���Y��EE��>��k£�\�t��,��Ni�,���
��1�@2�i����,0r�b���y���=ڀ�-9�l��C�� Y����ǻr��55z1��}d}6��,�w]�*eԕ�`��J�A'�P�V~��<%}���[6�ey�����)�Sޮ,�i�\����&I:]�"�ix����#���+fr�}&&�����>�RG�Q�/}�k<+O����1����"�#��ނ<ՌI(&
Q�F �FW��v���;*.Q�m�gg����sA��{�<뾎�defu�m��vs�ף��
0\s��E�ݼ�<�L+`�җO\�.t�S�|�K��]*ht��+5vsy5��H�.}(����=p���K~�-����zUyB�QF��o���Ds[��xtO������S���M`͈!ut��&ҳOQ��U��aj�����&Zn�:n�Ӝ�\�T')p������i&�����l�#���0F�������_Ab��/I�6���N�Nji�[�f\���󵈱t\�Dŋ����vk�<#�+���c��?L���h�4༔U�}�#���J��K�gfGÖ��Z*!,��"���"ixi��n��͐�#�IZN�9�鍠�;���J���
�aQ'Zk��ٳ�>���9\��\s[���k��b�vAҵ�t�k�X��$mg�b!sMͱN,Y]in��B�=Q^���wRZ�v$���f��3���R͔���[T�\D�y`%��[=a�C�y��-Z��(��( 6,�4It<�}�X�c�p���m�#m���3:���N�zhҮ���K�����w��|����o�h׈����þ�L��ڈzo�@��R��)F�:r�V�gj��T56�ZIo��d�v��x�Ӈu��!v�Ga<!�j��sȧ���XJ��,z��%�O� Jn��;.�v�V�'^�R~'~\wߺx�&�;�ټ"�{��O���(!G�T��No�7�1b��i�ʪ)��t氡t�:�q��S���a���Y���jxY��w��<�L%�%bӆ�z�A d�DL	P�b��>���a`�V,����D)��l�ԫ6�5��<D����z��X^�v�72��Hyy�y%K� �_��_s�9�t��Y�
��5���~QI*_	�ޖ�1�!P�o�A"|�����^�L�(��2�4^P�
H�V�߄ţ�w�q�`�i�'���5¾�.��PA��-�+LQæ�����U��n�:�m�ɗ���g���c���b�<���������M�Yt���ڳ��)Ŗ_G�$|I	|o�0Y����łFS2�D��DʃL�-�4�:�����'yr�'�H����)dL͈(Ar@'�G^.�Is�c6�7��\o�A@��}���G�t�sOJ�ګ��t`��Kg!V��◻F.�æ�7��璦-&eF�`uX,^��2���i�&��X�B�M�(�ح"����t�4Vո�#;ȁ�����zu�_����L�uk�4�M���7pVI�ɬ(��=F̒D>V����>|�# �`���������Ka,��υf�y-Uvd�w��x���U��.EbTt�M�8W�Y��75�+9+��URtE*uN�Ӛ�dgT��jx*0��B!a4���Y��~�xV��rw�X_9K�*��|�`�Ҡ�FN��qG�;j�z�ӝ��kN����;u�7��=��﮻&�3+�q���&8���k<�����LL�|I��^Id�FM�=���ק��[�����+��[��VLt�+s�%���T{{n<1ifcw�ZD�T���1��|�e�{�3j5u����E�Nχ�z��G��K�bt�ϼd
����:е� ���':����n<g=t dW]��qt=��
ά�ԗ�#�2HZ�㧳\T#*ʼ��x�拻[De��fuL�e�.�$��s�:E��}w�>{�3� ����)+"���{�پ��ؗ� Vt[�X�|Â�{�^�O��u�.�Q�9ڊ�����%J>߶�ED2�rZӁ�����s�)Q�*������S6�T�r�ڼ:|ni�.��ag=
HDtA�`�Y�Y��q^�6�	/�u^�����8zu槮tΖ
0�Y�x�ㆫ�>s��9ح����tj�9��=߁�����%B�TD�C�Y�3��k��'�U��F�jo���\4]��M>��oI�HXV��V��R�C8Pyl^!���`x'���O(���2&W�/��!�=��T��|<�Y��9�ʄ���-Թ&i�/�H�������No�lXG�GD���Y�t{��W;O��]8&*6���Ε4:�D�R橹�>,[�5	h��W��P��=��]w���)�ڒ:y(ߟC�������H�p`�'Q储�
��0�3H.n��4/i��N��Q����>��9d�S������EKѲ��j�@��j*]����D�������X��-��"����S��5�"}����,WSx�˷ªrax@�>'��vk�25�,Xܭ��};)���xc�9�R��I�k�ҏ8)�s�{������[3�dϥs�$��j���!��1�(����u�Xun�gO4��X��*�n�uc~=�� Gwm�ښ��]���}��'e?_��d��eWq^
�=>;�[ew�5���!���_���:Y��7�%0T�N�J�wrma�b^�����ޖi�{5\>��Y��a���&ܦF���T�
�9U,�۵�F�e��t౼­`����^B�*����L^,u���������)�T���.�֔b�Ea��s�ݛ��o�ip�:ENw����L �o�e]dib��
Q�1J��5;��\$��-(X?$�5	+���W�2;�����C0l�s����Q~��D/�Y���D3�%u��F����Ş�R���M�*h�i�A�sis.�}�	Wj��cMoB�s����{�}�~��ΗT�[�s�V@�֕�<v��EB��6<��sָqMΨ�]��Ƹ� ��ze0-����T�N�e�T�8R��Vhk�GgV5dJTF�XL�:� �<6�n2�{h�p ��؛�'c�Q��wi���6a�aC�*�ز�Ͳ2�����1u��Еm�E1������n�������?x>�K]��CU��	����\�Te��$G��oq��^����w15r%�鶄L��0@t�h�E�����yN|t{5�����[3p&ɻ��������Ԗ���o�=���o�~'֌��`{v�[m�m07��C��5`6R��Ӛы�<��𒎊��-�eLn,!S|��x+Ј 3���C���dQG�ͧ�|�����޼&8�yו�z"b$g�~�o��4Vv�=�ZP��u��^�褸i���^���K�EM2W��b����GEb���÷>���@�_+}��������J�����]8#T�>����vO}�KJ�J_�~&L�Z�h�d�%�P�W�}��x���+�i�Қi�j[�'�T��7�;7���K��?/x]��֔f�6����N�Ma�V"/缝�;�u���0Y�lSQѦqO������Y�{c���MUˮ�8���g=�T�w;��SVʩ�ھ����U~`���Y���Q�]J��_�Ly��0��3z.���t�U)�:n��6i�7v�V����W/�}���/v�����i�@Y����-��T�BB�#x�i���zτ��%��츞�C����JBw&�NF%Kf��2i�mH̿3:&Q��=H�{{�1����
{�a;�08o��wL�
v�&n7�����s�1�,g�_fŧE�X?�GK;n���_�^hi�Y��WU:�9��i��iI�0�j~��,5-٩hH߀
��G�MvtHf>L�
�ܲ��gG.���0h���nkDŞ�)H�ˬ����XAɱc�ݖQ{�hL��zw�x��j,��37d���1��20�q҇R$cXo���{j�]��[��T�F3���:�L��������6ѩ�B]f���si[%��y��m�c�U�X��K��&�{! �n�ֺ-PΪ`�G�U��xe�����ibÄ���~��� ���T�`�v��k�'dy������L[����NϚ��ODzAK�i>�+^|z�܋�dc�N�#����J�2y�̒4L�"$�)�#�����i10뛙!�'��L�����y���Bu�6 �`"&��ں��(o/̏K��t���a� �նD1a�B ]T K�4�0%��t՘1�q��)��(5tΙ�����l�9�i�i��80��f�w�&�#�{�^�C8G�W�.�c,������8Y
'W��u��X�ք�P���	�(��T8�-�%I,`���5�3�f�|�`�ao���N��IJ�2S/��M��Ȱ����j���rܵ�X���M�>쯳��xI_&�U��0�[�zENk�b����e#U�2�)M�6� ���η4t�*��Z[Z��,�lHF�RR�������v.n��p�z�ǧ:�g��|g⅃;o4���s'�5�Q�"c�H���`����qF���,.���tS�?��Ƀ���
�G��9�[O��ߩ*-�����O:[�X/B�O������{�z�ъ��-��c�s����fL����d�/T���}5�!i�v����Fc�U1̕P�cR�a�G�@��7��zY���Ƽ1tg����J���jD�#��KW+�8��3<�( �]K�gb"�@�!��_�{9x�6�ߗ����p��v���<�Mt���[�w|��c��i�>��$��G��D�y˖���n^Mbot�Ih���g�$}�F�އ(3E�!`�9�H�%Җ۸��YY�,(WWK��ExA7�x
�レ�!z�:'R�9̫���>�r�b���SV����%YU���3YBh��2��q�:�7c� +����O��rj�m��zt~=>o����1Ļ�+]ɳ�gܞy� ���$��ן�D�>{�}l3-��g%W��O��x�nI�S.�O��}�zMO6c�L���`΀ϭ���<�(�La����c�k�l���v�׾=r�Efd��}�R�!�3���|p��w�����:?w��]wɚ�*�gǔ�%�|H��ޥ��㞟:�;�Qs��SZX�g��"�]+�w��Z2Eg��$���%�]ȥ��+'+H���z+���0 =ϫ�^#F(|�L,�P�M�ysZ"K��{�;N��On�L3�sb��*9i��
��W7��[���=������]|՗T���tA~�o^�z5`Y؝~���2������ֳfj��=4�j�Qʙ�&n�d��l�r�#}��=�\�l��|y�r˦�h���Ϸ%����y������pu@�w��'w��go�xY��t��Ğ�������\+-����
+2\��AoB�ڽb\]����B��X�7y��T�$��ߤ�"���|��?-k��U�&�UXc=�խ��o-ف���s͕�78G���~��
�S�����zU<׹�9�ٻ��y�yk+Z�Ξ���1�Û��	�wF����� |�8x�U�H&�d�
���{��z&��ڒ
����\ƽ�ӽn�feD��uh�X�y��g;yMOp�U���w>��܊ٮ��=��oO�wt����i��}���b��~ď�Y`YǿV�X:�RA��N�d�P�j��ܜ�/Nv�B�Yد�M=ז�)!4���|�9�G�Qd���=��_z��Z�7���Q������-��wq_��\��z��8���p���d�z�������ʺc\t��c��ӒI���V朎�׾'������/0�z�p�z�a�Vٸ&��Zr0t!s.�UƊczn�_;�&q��mAB�������$v��mܞމ�h�M8��J��c�o_����}���u��g���H���4���f�"'#M5�;J�Zoh��%R���⩷B��:�\\�0�Ń�(^�Cº��k*��X9lI3&p��n��U��o\ˇ�D���F����ue
Y���틯�˿]�x�xv�1�s�o)t*��3��{���,c��3����g�,N�I���t1R�Gh����Ɋ��Iun�nȎ���m��RҤs-(�,��-�@AŹq3QW<�;��5G��q*�A�s�4�`�����#w/A98FN�r]�r�ԃ�]T�1]`JM�X,�3ˣI��X��#P�^Pqe��R]5�x���x�򻇩�8:ٍ��V���f�C�6� ��Sk��6��%#qR�P�vy��q�c[-�@�<�ڠ���@�|:��k9�sk��q��%��q�V�Z5U�,��q�V��[��@D0(TrC��7���M3�v�- ��:)���eԹ,k��jኼAn�lFٰ�6�m�
��H�6���D����Ҟ��{[�ӏ.ݼ��s��1���k�0�e�nw�nZ�:�%T����0
���� �ruٮɌQ�;�Y�W'X�V�����Q�QǓX�5��5�t�R����[��7�I[aT--�F a�x<b�;���:��C[��٫s�)��mnI�`�"��ѭQ��qy�g+n4��TA(����剨Xq���y�vꤱ�x��k�uY݃A�sTv�FU)
BY���۷��6���ht�WJ�Ԧ���[��j��n]�H\sU�I�`��V�İ�H��e�RV���i�$/�f�[��X��F�.h��o^nWrP8��Č9g[ �N}�D��5�KMum.��3Y��v��4u�ۍ����:)ø�#j���%�훈��K�b�j��-����M����C]t6�)����\���u$u+`Z�Ѹ�̅����d�D[F�u+��n�Wc�2��k���5>���D��\�ɁM��Bqs��lvb��X�]����A�ɢ�[Z��V�imG�{��Gcq�.��@�j�rp<��ڥ�۞خ݈��w+���!���\:�%�D��k�p1�"��DD�����(i�?�2�~���e������\��7�߳����lߝ��|a��$�s�FUN�W��uc}���Ś����a�-8?/���H)�
΃s�<�{�{��qFz��^B��I���aֳ�+��g�d��_EY���9�,��
���:����r�ޚS�hA���O���k����M��ͱ��',^�V�V�}�o|����o|�@ά{�tC�w�7�ߺ�&�޴DF*����B�v�6���j\�a+[B��g��)������W;��&���׼�nZW<�Ӧ�7UiֻZU[�*�]�HW����"нF\��oJ���<�dv�š�K�C�*a*�u�q"}�o�W��j>���C<o�B�Y��n+��}�Q�����c5_�j߃T��5�ŀ���a��:���$i啜\��`�ݣ0$����N���b���[�#�U�GgI���T��Qn�U�9먭���bn$ћ�%��"�}ڼI����u�Z����Vvz|����c9�+�t4�ٌ�A��[�{�'l]����,i\f ��nH����{p�{z$�A�Q�Y�޺]|���9繙��X�uw�:5��S�9�JM�ے�:f�����[f���W�q.�%��yq9SǴ<�Ļc�b�17u��L��u�B��hk����Y�r����z�[x��_4ɹ��o'oJ��N����<�F��I0W�֍\����n�=����Ѷ\Wb�˛*Z����Mj`���*��p�ܸ�1E�L�譣I�V���z��7�Q���	�9������+uy���y�����4�D˭�G[�+DE�Ь��eŪPd��8���v B��#�2��Ƹ�ں4�Q3ړ� Z�RV�ie0;T��ݱTX�ki�*��Qn���8��<c��}�A5^Z{�o��T��w�vn)Y��=���Z�=mŏ������Q������N���˼r����=蚌��i��M4�';��x��lT���f�uj)X[���KKh*O$�Ӿ�7tѭк:9N�� Y��A�:l���u�4,/��B�ų
@=�dfo<��Vx�8ﮦ���
��M6ńt���^T�/�<@'�O�I_'�3$q�����D$8�d_wS_��U�� (�F���/x��U*��i�T���|�.�}��|�J��/LKN���x�'��}(�:%��4�y�5��t���>_gNb&��������r��WK:p����T��~�O�
 �=7�u>�A�`��D�l�t���e|n}o\��$��vs}��K����y�krx,>2����1']_g>�7�V;Q6K	���T)��V���eį�r�J����g#U�｜pg��;5��R�3�=;%��/\O�f2�k:]��|��J|D�)If���O��U�jV)2�*��}����v�i�N�ͩ����PeM��*�l6������*�,����a�${HO�}qv ��b"�MG��j=�,_��j29���U"'���!�P�tf���i[�'��ƌ�=���#o��cH�V��v�D1#������6�P;3?$�K�d1*�]V�q}g�;�C���N>eZFz"��@E�1��~i�f�bꑸޘ��|����Vt��V"���E* Պ���������,XZ;G1})��l�J�7{��b�BU\@���d�5��i�v��Mŝ$�°�"�E�B�{�^�&�����ֳZ���xs�"�psٓ��D�
-���J��a.�_b�"���ʆ�|��ӧ�������S:�"J�9�ּ�!�bf3XXM+�U���n;�a���\���g���\���\F�|�����;�x�,��u=2z�� �|,4ӣ�9�
��'���%:N�$�n��ذᕼ�xw�Qi	 |GO�7��\��~��qh���b����"�H �S#W�G�P���c�庼Xg��X��1V�[.����fH�!GZ�"f<�� ��{��xXuQ qg�EA�G�"���v`��GH�>i�rorc�Z���d���۾V�����rY����;�E�D�BN�kVk��E�9����r49jIW{yM�c�8�%�r�B�ƚ�W5���|8����maF�W3��/���9�r�[�� �K<:>����	��ｓqF��}�XQ�/:<9�P��ِ����R�#��#��S2&M40)�/
:/���KE��B�B! $
���϶��k\��y��:�H�'������V��f��W�ڸ�	x]�v���l7]��Y���������8�=�}��Jji���t�s���\��މ�g��s��ZGvl����y�:)�:iә�|{2>?>Ӆ1@���	J$$�L��"ȣ���K��^ ��N�}�d���8p�$�˕����U^QQ!���zC��B�
uLd��ipѼ˛��f��̫˭�B�hB!����^w�c�7�}��O�d|�z�x,bjtխ,��/(� >b�w��|F��渲$���W8���z���קP�EVX˙��N�t����F!���?��T�CT�����"0���"������f�g��$��B��r�~�0��C�f_�Q��K���j���o�xXl�4�]T3ڇ{�x2oP9�0j�����4,
���K��Z=��~��	0�	�nk�
e���+׺�dp{�KɁ�~G�}����{긡tL��U`��<��]_���\d&vitQ�p.8n�f��VË����\f,�g�� ��;��^c���U7�Q��n��f�ᄉ�sKјQ�r�?DǗ�0x��i�k�u߅^���e�i�D��f[��&�>(�e\_�U�	J��_��T�B����;��'O���R��$W�"�V�����R؊��U���c�;8��L�Н�w�[�W�/��B��g=�׋4�e{�yZ
8&fd��.��R��	n���g�]P������p��yJ�|a�nq^3�ߢ<�B!a�z�^1=羟;"\j՚f�^M��M`Μ/=
��(@ć���`���.^�T��8i7�w�R:p/$�-5�F�<j&AaM\^Q����5������#gL�mL"'s�s��zHO�i5��g�>�Hrx�~����iAGt=�����[�vz8��W�e���s7g[��u5�l���Ѫ����[E�Ӎ,r�[պ�9����ɹŮzK��r�WC`����ݴ�v�
�\���oI�����A<v�CxǷ�]W��Yۦ����mv�u��$p�3t4����L�^�\�Ū;x�vԽ0���"[،ts�9����Vw@>��kuO.Ӽ��9��u=�ݹd��ݔSx�t��˒�O�Wr�=��|{x������~�]p~r	�:�m�����di��s�[��a!Y�.&��_wxp��z�[m�R�rUS�\#�1WE��z�*�t�v�o����@l����G�7�V`ߍ��TӡSLsM�pVa�U�ɞ��zD!ex���7�LӃ��)�H�/��Y��$�@ o�z~&���j�U�]��zaz��v���D1w��k:�z���'b�I8o��t�_އT�D�S(�O�<���T�$x[���{ʾ0��W��m��  �,�T���.h�ɏ�+���`��f��cX+:���حigEg�A �����>�Ԥ�w�����s���E&�,�q��i�&�9եΫvdlt��'�]V�7N�y��5�,K.�y�o��8Y���̰XQ�嶹ụ�oޥ�nV�'w��Qs����~I}(@�P ��N�����v�E��/I�I�Sr[�]:�5/�?�7"߽$aʈ�j��G:9�'ā����2g����2�S�Փ${�G�dLD���CH֑q��cd��g՗�̸|m{�ly�s�_�ɲ5\�ՍlB�+�c�������Ssx"��V{6�2e�w�{��E��ݾVʑ��b�����,���k^�D\��[jK#�r8���H$Ax����l6�����T��߅�7��{�-,È[�^��O��*J�+�Oz�JH�}��U���2Q��[Z���$�V��9�J����Y�7����S��X1t����x*"}��9�!rs�y>8V�����X�m�Ny�mwiɹ6&��BR�Ĩ! �K��"O;����I�!�f5:L�g��tm�Xf��j�h�%v�Nx�y��K��[��f��æͫ�pC��Sښu-�=2/2�����p����0�G	;��v�����᧽U�=�L��J�N���gWd8m��Sf�}��	i�޿�]�d�ʜ�y~k�6Q�{8��;�eg��a 	 P0���ǵJ2�D!(�b���\�j��4_;y/����R��~���k�Zlwk��"�ʌ4�0�"��a�����|�|`�uOԯ�����@h�9ζ6���g�M���TӞq��oX�����x�qzZw��W��ç�����b�-�����Ҧ��Nc��H��O�O�U���g�b�F�d&)P�
ĩ1"P�I��(�J�(�!����x�i�~�������&�ӄa�B�B����k��1�I��#i�T��XC���SSܟ��(�1T�BF��Ѕ�q��g��O��N�{6�a��߲Oz�۬�t���i	\ʳ���0yz��jM�A�F�m�`@#��C��w��[���q4ۿ¢��ɬ��/��q'Eg�r�_�P��ꘙ��7�f��b�M�.X�9M�nVњ=�W|���t@!Y�*��;k	�'���J�יMa�B^D�4��^��-��˝`��~:�ݷ�b}�ef���$ @}2��щ����4ષ=7�:a�VI­�Jj�ҙ�m�(]�$��XOM�����I����f�6D�wdI�� %�ۗC�C�,�b	&h�dǉ����bD�JN�u�a)�iGX�\��Q1����7��ܧU-Wd\�YS"�I���Uu֣�FV���o��|�y��u��g9�z�|<@Ӎ����W�d�5�'u��D�E&B����wf�YWM�������`�5Y\2�k���O��T*$A>��о"�Ƨ�_�B{��TȰ}e��pH�{�#hA�,laSb[���A��Ut�[sci��͝y���p�4}}�޶9�����h�8-�������3y5�H��O�-�!=+�N�s�t�F��U*���8!s��N����ɷ�����%*HA�z����~�v�5��$�'���B�h]��<b��uꙒ-ұ������p���u���>[WX��O�O�:)KO�����҅�����#80�;<`$�:�@�@�>�IxH�.�s���׆}����ox�&a��f���.��/B @ ]缟���w�CݯZ�j;6.e���tJ��&��gH�����}�e�ӓ'��
dG/Q�|$q�Y�>���Ԉ�+S,�^��aN1�wZ��J�AX��/*�0~���hUS%gj8%�&%B��{7����|Hj�d��1ba�ѴZM�;ŞkS�����+4�J)�bF�L�f��S�p�Z]-�B�UlHX���t�c"���m�%�.n;>�/nl4����;#1�vb�ۮ٧����B������\�]�۰sm��ԄH��k���&�Er�ؗ����kt�&��In�jV�&�[Kb��PWUDڃ���ѵ�m.�ʶu����a�f�{u\s7i܋�v���>�6�k>p��bz�;9z�&%2�ú�7���xm�J�_�˘n ��֮Y6r!mCnvm�X��K�h�#��5�0@b���p�}��y���MWt�4�v���t���4扚p;U�&�D����W���F�s%���HIL��$""dsPB5
6������F f�������+(����zA�Y�2����	O�𴌕�d����R%� _G�e�Ô�4����4^z(�)B@t�d��ǋr�\'��/�������.�L⮌|�W２�P ��'�쫆x�b�^����,�yz^	��]�I�!�$Y;�w��~:&���g5-SV�kׂO��yK"�~��B	�7��G
Fo�X3����gJ�����5���Lݠ4��I�ݝŇ������f�Էpn ���|x<x��y�~��`�]��4꟥�:F^�>��7�oSXGN
�}¯�$�Ù�zixү�׀�igk��誚�t�6�]5|�L�p���D
�ڈ��v���� �%D����`�d���Kkn�P�"6�8@�����
�<����fSw�]G��MZtB3�[*�1��y�:�a���1�7��Q�C#^ Fv{j�b/X�yE:u���B���$��,â��:_Ef�㹶���@�,�����!�O�����uu�
�9�]4@���K�Ί��_}^�H�
>3�|_=+�>(��8WBy�2�e˵�����p��谓�o�4����]����2��x�a+�/*@����zpӇ��)�r��۩��uL\�p��n��Q�]R(y�����8-����L8^]�0�:G]��~�~�x|��etf��i�v�8��Wu��f˱Z�R�kS}����U\�D��FbUi�V��OЧ&3t��fw%�&S�������@����/�������T����)`�t�Y�^�r(]���+�ɚ���L>�
�d�]eb4��$�0@��*���)�	`�e����>����&d�IZG-�L�;�.*�#bN�*$퍷4�S�H8d�i*n\�"�ɑ����gOR��V�G9��zpT��g�r�� �~s�.�S��t���l5��}�w�%��n��=�!{�Z�)�������nn��i���T)0��-j���`�se����msڃ0���ٮ��M#��P���' �(�<����;����{}ˎ��u�G���@#�{%c�\央/�`��hI43'�m�6����K�o��4|�LG	3�{hdL�ץ8�Θm�\7b݉���|��]�㦡��~��=�g,��^n�=�ub]�omlt�9|ے���ؠ��Ȼ�R���"?�a�E%^�1$�6��V)^��N��<��Qu{Ƕ.��s��P�bJ�D]�>�a��p��w�)t�51r�3�"�V:�X0�mv�&��LO�g@�=�5+��b�ԡ��z�cb�ag�H��4O]k�[�����^_�b����j���h��qm6�ulZ��-�.����1���DDj�vi�>�z��u�i���S����n�����թճGx�s�l�X"�=�_�\>�Y�<��$\�`8��n��p�������R��m����7.�!�rȝ�O1�]U_7C4MPX6*�����GN��;��X����37b�c:��-�����A� ��8z1����[���~���N�Wz�/d6}7.����Lv�gg�@qg�V78q�J����e�*��Q�OM�ב~Q\��{���|���|�RUB�{͝���-�'��f\:b�Ul�aw�I@����<�8��j�06m����}��^�D=P+���������W[�j�3�^Bګ��bqe������xޝ��yk2:�<�b�-�{�}� j����V�{=��<�oy�Wl[�W�ۼ#)]��̶��g=�	c���L�uM��6e�uk���W��*U�CT�s�Bn�>�����\��N��c��?]K������_I����T���Cϳ�h,��u�;|^C�W��*^�|�*�!�i�7���F�3�՚��������h���9�M>>�V��x���{
��\������?8���N܉�(Z��kp��ܠj)��|�t��#��UQ�
�x.[46�F���^��Ay���>�Vv��ט��ˎ�lO^T���Dqp[W�/d>���7=���:*c�A�-i����^��UL��c���m��x�jR����Z^��ߔ��0��:^tq��9�[�lu�`faW7J������[.,n��1��Zc��'z�U�.�)�����S�"�5z�N&oHh�b�7P"v�wYq�Gv�`��.u����q�w�yr;ˏ����������&S������ݜ���Uc�O25}���b�sۅ��|����)&{��{�����i J��n�_~ai
��( �V6E�t)��
9��E�}�N�"�ܺ�J5,�ao�ۯ�q�[9�~�#{~?o�{<;���"�2U5�rc/zM��!f�a�-߼u��s�q�[0,h�F&sc�Taj�\�4�DIA>3@����3D��Q�F�ڛ����Uԝ&Cyk'o'j���|t��J9m�d�+"�wf�L&~ڙUK���ܩR�f���'�_�H!HA����LӇ��r,}�^`��/���� ��~qⅨ�w��&�r�*�i�l��p_�3�,(�M��  ���򸣢f��FGM׺���8o�r|^�Rƿ̬4��k��Mv�eXX1-����FUм\g5ټ�f�����8�����5���K������*o��x*:/����-��������KEdpǾ�f�%v�s*fYRtH�j��Ogb�m��|�ę	��vW���voD�ۯ9XGE�f^K÷�(�X@��pU�����8�aj�=.�ӳ�o�N���8Ws��[3�^����f����7ёژ��rEH���2ۥx+;�^� ! N_��^#N[�:��/�}�.�P�2�2��G�3 o!b�f�����؏z
#�'"�{�-�R�"c�b׼�
�Ʈ���*ӈ��͡��Q����bw{���������C�RT�H�����V�eR�yQ6�f�Z1��? �@]��ϋ�P�4ۑd�e�ML�EM&��d�X�����Ί���T "���f��
���DΜ;Sx�`��E�o�C�|�R�M$VH�SnRp�:`q���4�,θ��/=K�uv���r� ��*��%L)Q
¿��Ej�_|���:����}�ٕ<�U�f`�M4��u��DOO���c��T�2r�7���'��= $$F
D�8x���Ysχb�'�+L4p�k�Y/�I	 �w����O����BY\�ν����kt�:��\���%�$#ҳe{�t�P��=W�s}>8>�	˶i��Z��� ��/���!�a�~�K�K<.W}��"�'�����&4"!/gު^(Ӈ����U0�j��MSj�*p\0���OD"&@B;�y>�V�2|]��g�0�X���;�N��9�0눠���R��l1�U������<(���� '��veI�q5�;�*].���P���E{5���M2�i|4��ۥ9
T/^�f���������wb�;OC�_�N:�j��89^�3$q��\Q�v�v��m����X9��a���^=�kl��b��S�]infnt���K����D�-�b�Fx#�����;O��ι�z�x�W:��Z�pm<�;�#�;xR�Z#5��#����Ҙ�j��0�[slIu��Sm�#wHø9焀��;󬞚Ћݪ�s^�3Ƕ��c\C�.I�i�zt˳Gg��~�U�V9<0����c��ݒ��ҥ"�!Y��,�qn���a6ZU�{9Q�I��{���x8�:��m��ҥD�NJ���ȃ�/i�ɭVE����>�G�@@�sҨӧ��ZY�����kv�l���z�����~t�>W�/%" G�?����
ŝ�/&����/*�.g��hP )#/}]�r��3\�zc��_��P)����ek��H hB �7��y;��O��~t�$];��MYV�DK����w�Σ��Q ��k�N��ਆn�5ZјO�OD@ }+�������;�_ޱ�F���W=�+{��*:gҼ�= #eH�;U#yn-7��f�E�{n8��h����W�Kq�a��n��kR�lq�����Z�׳����	�3-�}oT���Uu�u���EdX����J:pOq\I�p]̚��G� BD*�+���Tiè^Gԕ-�n�m�,#����C�\'Ո+������ @�%C��G��D���"�d#'���Uv�ڢ�4��S�W����jk��j7�����H�����:&�V$������� �F���`��O�x��/FVf�Ja�&a�E��	 �}%��-Α���6WS�Y�I�ubF�c�r|t_u=��*)�Rʚ&[��Y𨓾ɮ�a90�r��;�Q��BV����r/���^�����<�vˡoH�].U������q�P	t��.^ʑ.~�\�
0��ϸ�%6���@�$X-��iB�|z�(��M�|��9���kQ��vw���)+�L ;]�+�F�u�k��	��+�k���K|羨�,*%:��=�ꎭ��M��Z�sb�m	@f�ۛ�%Ϝ��u�֗L��Ŭ��=��zvN�{ܛ�w���7�xQEN���@�"��Z褙]Q�!��Ր�wiDL)����6�/
:+g-�{��QiH�\�;�=��zT�1c�t����o{� |	����G|~J�ӗ2�S`6괡i��+�o'���q��z���{k�c���eq��ҋ���q!J�&�{
ؙ�囘(24�Q �뺌Z;��A�8�`�;#K�[G��xq��F���Y�#���&�;f���_,?1��'yh;�b���ml�>y�	���<�E�3�[���g� H!�x.V�+��,"c��zg3�R��GD�*LD�֒P�|�k �A  c���������O�yWӥ�.
^�(X}�Djp����<_��>���j�*eԷ2r,#�>k.�rx`��B_*r��DR_s���C��N�)�|��{�P��;�]���%t�����i�2Yvv ���c��M]�h1Q�y���LG/���?8ٟ߯w<z^��'uf��9vng|��6=�]�±h�pz*0��kQ�w���ADEIَ/���Q�O���(��@��S4��&�|N�5^�䖪! �p����-xf�.�/�pΉ�{�/��w���R��s�s~�5�ua�j���)taK���GO�����C�㐤�
 l���׆-,�ܿ+�GF��Kw��	fr�i>���G��g� �����W��{j��oҾ�OEf%�Q�Q�g�K�+��� %2��҄�HCl�I M�Ljv/zÕy�ha���|�X��|3&������B��֥[E��[2/�sP�B\{I��^��{ ^Y�9�=܉���0!:F�v����XB]��'N ���\3��6��h�}�$�D��B2�n�?w��&���1���cu�׆:.VJ�"��ס8���B��p�>{��Zѕ�f���(�~P��{>Lb�"�ysvt�a1�B1Ǝodh���;���`IY�)χz��/s���z�۩��P�.��~�^��8mo�Y3,O���<���	 ��h�^�Ƴ�b�M��>�*��i�S&]5}4�����E��Ĥ�	@pҲW޿u\I��eg�k
�	�}8�;C��I%P��wsZzEJd�UMMP�F�#���Ⲿ�b�].rX��t*H 0�>�|]�E�?y5�gNoqVӪ�IrԹc�7�N�B�@#E�s��*p��Z�:p��9�>P�)�#>����4\<R&K�OA9uR��6�1Wf��ۿ�I=�e����3N����4I��F��4��x\��c	>Wl�s.B�x*A�b��:Y^Gu�[�(d&B������}̥
E�Y�q(V.?R���f'���n�M�Hy��,YM
/�"#�\���=�0F��>��s[9�Π��S�n�'V|xj0<�9޲�7G!c�6��M.�Mcw87^���yū��D��j��-�+�1��KĨ9Y��4��n%���&�,sq	�L$@.v��Ǎ�3�b���MF;;�\i�7[�#�o	��<)؊�����n���j�
۶�p�i���!����\z��!SB�H�ie�ڐD\d�ƭ��$l����=�g��	^;jg^7�٦$�J�`�#�5��XeQ�lô���f=&��7ۃ�<����{�wb�M�4nVw�ņ��,�t�\�����g����+�y�@����F�'����Ƿ��ͳi����<���vG�y��]y'� �	9�N�������ǫ*9��MqYGB| ��A��%�:/R<�'Ԧd��!ҿ����ϭ����}��./D/B�@�ޯL�i������N�0/�ɢV"JcAU5҅߼��!�K~�)ߥ3rz/�~�����?m��<�G� BI9�y�$�����*er[�@�Fܚ� ����T+8p��R��@�
1=�웆x�վ��\������酝>�{�}���my����"�l�m��mL��6͸b�v+f�j߫���px�����,uN�o&4�����F���~�X1|X�y�¼�� �-�t��9ӂ�şͅSNj[L)���T��(���/�*h�YcF�zclEUb�B��fc$2=�;���c$
���{X*}�H���yz�,P�'.=�����n|��T}zb�F�"Vȹ���W��N�����Ľ�ӼrF�kb���t�&c+m7�G��|)
k��%�g$����~���K�}�D$9<,�zD�>{�(얱.R~$Z2}y��TC7��\�l�B]U �k��ܛI�}+��D�#'���k��
�U�xL}��=`Hp��9��J�/e�<�Y����a���i-��>���+#�޳̧R'*��r�[�aGN	�s�������K�*(��(Z�go�O³[��~9�{�����R���]	kL������vj��z�/(.w�wj�U��s���~x��w�}�{]��\�eg^�}��׮��,8N�q_��R%gn�_=> !/4y1{�}7�E�O��إҚ���n�������y*�p�;5�^�]4��={OJ0V-�-�'�'���������[�m�
�^�����]r3��yD_�:>�cGeNZ�wS�ȏq���'�Gj���56�������z��b��xq��A�|q���?2OZv@�s(���+�`��ۛ,29�\��po����������gj~�\����6e�0������� HF
��](]#�u<"����oZ���Ar4�D���'�-I�@t\�7���E��p�Ҏ�F�ŷ4Ȃ�{��2����2�3K�~2��E5Q2䒛���蹲�����فD?]{�9�Q�k�r`ы���ѝ�}�J�r���j��n�vu��6R��Ы��..��5s��v� ���?�x����S��-�|P�f����:|G�Q���`����������E�eo�5��ϯ��& @��23H�ܰ�+���IQ�
���y��8h�=n�]$],u������<����d�����W2�Z��X�D���=��L��̧ҏ/1%�T�(�[�]_�,�����y%���\t�L�
niӫ��sТW�ȑAߧ���s�T�;S�
�,���*�A�<����]����V���(��8[�tK1=�<�ܨ��ò���Ps��Ƅ�`i @��8��&}�yc�uY���\Ø��dA�������:nMA�.c��n�yy�iՊ:��6��r��M��!����\�o�S��۶�K�"B�fp�F-2$��BFШ��B���Q�7&;{���M^I|�J�����#��'��u��Z�)��3R�v{���=��)�L���s��;���Fɬ�m�h�g��z�)خ,nM߰�����&Ź�mT�UNo�d3��`ΟrU�s���}��tY[�kбI �e%��2+|�Wϐ��J���@�RTJ�3*&�{�ы����|A�7�+��GO�S:���}��g���ɞ�j�je�&����ߚa:��ꯀ=��I$�����}ݿ�|7���|�-(�h[��>�W���	��5�������~�1;Sz�c��z��!�/��l�*M3Ȗ�ۤ�M�U3��W2�z��yZE{ݝ�����G�7YM�t�ߚ&\�(ډ�t�'b�댝nDN7U.2�ADa�#a�koú,n.�J���o�(罗��r����_��y^�n�0Չc³��Y����mb�a~;��	�v���S�6��U���뻩���Li)��P]<3��%|�P���T4������U�ջìA�%n1Nȇ9=�zc��ȨOT�:Q�3��K���dL�ݙ�ϔ�7f�Ha��ߍ<�I���Z���%�X��T�Il�x�Q�o���-�M���xl�y�0���n\�X[Ï�_	��H�����;� &�/���ȧ}�y+,����yѷ���Q���r�����vB���ݻ�Ћ�k��{�ҊC���p^��9#�K��eb�ˌ��m@qS͊�V^:!�kӐ͌Z�N`F�H��	�J-D)��W�]<�e\�0n w	g��fA��k���'�,t%}����_|���1|��5�ۿ|�w�w�E��f�ȇN��:vZ����WE�o�/���,�`�}�grƽzW��q�n�n��E�U���7���عޯ�/�/8������y	�NNX���b$PN��Y�%F�5����/�W��v͛�����C������nTƩHa�ۊ�_:s�|{���٘
\��d��0z$\7�w=���~�s�a�5Hg��b��}�_��y����1oE�Z���+z��͈��5Ki��u��$%U���c�a��ʟ���53�t�&�V���Z��X�e����mརdn�i�����pW����Css�o��1u�W&���)�7��ֆ�bj�'��,	i��pZ�b�:�sy��4��bŶ�sj��^8��bF7�`����_��8
g�<_9�`J���K����Y����Xp�  �u"n۬讻Q���ݻ;k���@t��%�Ϡ�qWZ�QZ�al!m���VU8v:�M�ͷc�=��\���2
j�fn֮�,��:���v܂Z,�4�ˎ�7 �.B���ά�msbp
��F�%����\u���������b�%��7��έw1�qq�<�x�����GZ�#��
�ef+��Ma��7+n��R�і�)e���u�lpQ��g��r�2L�˨�ź�N3�Kc�GMvYf���̬��u���l�v�x�F��u�F��[V��n-�!�p�&�\�q� ����Yo1�cb�b�VՁ]-�y���̋oN|��p,�����[�v�ᄵ'�rT���3%���e�g:��f,��s[3nx�����J�4��vԄ�U��-I�-�Ժ����>�e�x!;��,��(������۴�&��K����{q�jL�j�4�[�Ŭf
��������8"�ON�kn�p�X��p�
LG#Z.�B��+�����06��[�5b:��q(��i
릅�K�3A��,ZʗfY� �]�� ���c��n��Ć��ËVe��L�%,�5�[�,K���ѥs��Z���lQ���8�����i����5�Ɩ|r�3э�+.Nn7ZF�)����0�m�+[fU�m��R��K@���R����o@�7�v�>���!�j4@Hcl�v�����ls�t�F֑��m�̰���+���F���tK�ґ��җ��8�{Yg��������3j̣R1����:f��j+�.�s��`�D��m�^ 86e�-X�QӲ����� �f32�-�\� &b������[kV�� �-�B�Ye�v E+R��sÛZ!p%&�� �6��	[0<�`�������zaL�K�`�m5�46��[i]*�,�:�٭u��Ҭ7��]rE�����u��~o�����c��GS˄̣q?ýw��]=��,�B�<�r.Β�=:�,n7�z�:&z��?n?/��ks�Sv%��uw���{v�����C����I�{����ιH�����|�����=�;�z	�j����mQ��L�{��b�~'�9z��]V+:�ګ�3D�s�+�J�6s��cx�R~����#mHS卞��̊;gU8$E�*���l�2zl�����ﳺ�c�Ԡf�����k������c���$�*��3��_kZ�	��ݧ9�8؅	T�=����{`K�0m�C�>���R���j�	<��߫��.�ÿP��{�[,�'f
����7�|o_y�L0�}�{�����g=u��ѡ��8Kp���si�h�{ÉP�mThR�R���D3P��{�df�*j��^j�t�a��a����C��P=�n��y"�C;셈MYY�a�:P�B��Ю��D\L�3����{�t���Q���V̭+��pƳ37Ӵ-%1E���yr��n���y��l��1�{��6n�/�'�Lɟo��q	��^;�LJ�-�ss�. f���|�5(�ꙮŶD<�2��9������U�#v�3�wӟ��S�N5�Z�'M��,er�vr�(儖��["�,Z}{R�<�j�ώ��<+����{��t���ó-�K�q\�[
Jʙ�eJ,xJ�jV��[�MJ��-��u�QЄ�EK�]��Z��g�/Y(݁��ݬ�%�㷒�^�7��Q�b�\���`�M�d�L;����k��ָ��:����u�d=r�)�Zg1�tֺ�H�n#���[�i����Ld̵n�Kb��w��[\󃌁�u���d�f]��ei���!\I�ѺH:4]9�ˑ;��<���f��]HKkSM<)�~D\�n��ɯ='d�X�n,��B����淳Q'cQG���XG�-KA:�K$�ph���k���x��G��qU���l����	�z-R
��Ș$Ľ�ʗ=��p��[W-�π_O�����|��~�Rغ댶�쏛���<>���=!�x�}if��M��ϗOTgm'�����=�h��
��ꛯ_��������=�_����|ӫ��|WN����<��qj��*���Ȧ]5��z#&�w��W��G�͜�S{E��v���4B ��~^��Ǻq�����%�o9[Y�N�w���^�#.~<�z�}Yš�w)��}{9?2|��c5��Vjr���u�hڤ��F���ŵA��F{'=��&�7mﴩ5	a�$b���W�W��_x]����u�E�� @D����'���r?zBD�RTL����v��� �Ȋ�D
�=q���y�Qr;B�'ڪ �dI}ԁO��j5x\ �<�ז+zPg�}fdsm�&�Mَ+����뛗�1�L^jt%pv��֧���2�>>����Ċ�	�4�Э�q�$�)"I��v���S�5�ڝ���x�A ����/��lr��]-��{�Ƕm�:���W[�G�^ӧ/��w���M��sݦ��Э��������@H��=]���;������9sߩ�%���%���tu#�\@PA�O�J/����z� ��xϾ��^d�w���OK�/��~�8>��Hʘ��e%�q�J�k!�T4Mu��b!B�<��vr���=0�b*I����M.������lw^�{[j�BW��B�}�^�x��=�''x�)Ț�eSt�d�/o5o7�� @�@%�w�{.����_����Ǔ�J=� �Uγ��Q���J��LL�Fm���:�l�G�z��UH�@�n|�|c+默��iOl����!RA��VP q��0ލ��C�}܄�Db�@��nE^����9Ғok)X�B�F(Y^��/%�[���3U��+rgm��.�V��0��,W4n<��  9	$j�s��e��/h�t舘��ls)�)��+������Ȉs���k���/7�t�u�/��/(�Ge������s��d��-���m�=χ�s���D�"A~�F͛˽�r��s������?s�[�~��!��*���#��'^���gU՗%��5�5� �9��NP�}K�g�"f*e}�|��P�:�x�6N���|�!�7��_�>Y�sd��MQM:u#ms�]�uxw��䨄"o�[�O�y�O�w�æ� @�R^$��w�'�N�e��S��>�~x�qv�l��;5��@B�s|�9���~��<���qN�f��e�Yy��" �/|z���ߡ�ֺp������Y��E(@א,���ϡyD�"eE�&����II�_R�1�Zc]�R�]*��j�<�뎡i
O�.e�V�j�Š��{}p{�K �!�H2hd ��S6{s�g�����-��7�/��h�(��䰃��Hv�t=��ߗ�P�Z��S�4�H�I$�&��7b[��(��0�����nv�Ϫ{����9���= @���]���?}i�uL:���;��:bDܻ���p��Il�ؗZԮ܈C1u��WUս����~dC��vu�m��Z�[*���{��3k>�׳��2��ݹ~��j8L Q��־�cH�L�B! fHS�퍘ny��@�]_|~��[[�u�7�;�P�6�.{�s�DMT�H��u鈘�'�j����Ɲ�y��Ο��}U�{�b��̕���$�0��t�_<�1$�^$&w>�N��|�U��}\���(�)(;�{�������X�M7ULuN�Oi����p=	z"���m�/�9M�8N6>6v|���@�����vw�g���"\�l֬#Ȉ5����/a�Gǧ��m�d���`���};q��Ck��R%�!!LG�)Bf|ݱ�<�Y�s-��w�R�:�cu�����:�u�۷*^��z��	��&q)�M�C����n ���Yk��W|�g�Z�͒ h���[bhغ$�ne^,ux�^X�g�T�Җ�5f�z�v�tN��];F5(:�N��\��Gd��5�ik{n�Ƞv�(�V�MFZ�nZ�gR�,�	ͥ��/k�F�/�4���\���RQQ}g>��p���}���{DY���GA�wO�ҝ#|77��iM��3�y�w��<�y���&�s1*�<+6�1u�#@�d�n��/A���n#���~�x8=_}�9��ݴJ�1*V�j���s��$l�2�V�p��E� ���ok���g_��t�rZuR�sC����m����(�$K����m}���|��>f�����<O�����̹��Ni�M�������[8��o&�_�z��꟢y��5��q�r�ӋA.ܮm�����[�X��=�߻�����~{���՗��Bز̂ ��gV=g�eg�h��s5L�m��_w~5�W��� #�g���Q��F�%�<�w�~�Y�)���*�#5��d�X�WX�M�Y3�,�q��s�Ύ�ww�pn���1�BFf%L�˨��ֶ6\�s��ԩ�}{x��~�o��x�5L���S�*et��
'z;!��[�f�*�V��0�@e|k$�JiϠ��|�d���>�}d�O������L���D��R��D������iu1����<�X���"�����^�����Gv�H�p��i��$%�^^���A 
���t�m��7���;���@ �%О�沨�Ӥ�M���Z�L����roowO��� @	-	�|�����߼��:���4!�sT�9���� ���>���h����k-��'�}�|>8M�}�̎��w�G�G�!P�USu���gϵ���?�Ds��[YK����ͽ��;C�ւ��&`������^\�(0��&�yp͵F��Fq\L��=����\pxDn�|&j�L�T��37��wιf�2�joggna��Z�m�w���^�]���.UQQM����}��2��%�|7������>���YQ��Z��|8��B8���g���fٗ.��f�?Cf�Nӣ���x{��)!ڮ�wwK�����>�����(������\��z��ϫ�u	#eG:����-m��p���w`=^�u�f���br?�^OaZ��s�c���xuavnA&l�WO�q����q�1��QU+o�2I� ��ʹ���_����l`)JDyD̞�t��{<��y��:��_}��gy�N����ر �G�>�/M��~$�T\��6ׯ�_��}\�D/+|���}��O�Nbnm1?@/��T�0f%dε4^$p˛s���cA;n�Qk����:��s�:�;K�՚��S�����޽�M㨗:��6Z�{�0�)/��W�7�V��$�W)&�[MOk�go,/23�z� By��������Q�]���v��z���Q ����3�U^jI8���g~�=�Z�X�g��0�����U�\w������EJ�!�L��?��J��|��[�>w{x�����Ϸ�bd�`�%E�r��D{���۫>g��\0\\�!X�� v�k��BN��H�R��෧"6k%ӕ�Xqu��tr����`�t�O;��x�57�[*��A��,�GC��UP���0��I�S�d�TÑ���r���,��!}�u��>��$�M�˗N��n��;��F7y�xO��� �������}GK�%������w�
��K4ԑUBc�V�i�)p�.��.���<n�\궼W~�^'
r���-��tb-�\�����t���ξ��n���G�`�0�RG�}���u�����+EFL�(��Z��W&a���/�o�ӯ��[��~]��{�J��B>?�o�zc�pF�h9g���	��jqV]ov/(�B�'����em���}}��[��M7.�*jJsN��y�����o����� �2���{��$� ���*߹�n�+�J�rӒ�C�[9h��;=��� ����j�+w�Wn-�	����7��{ ���bx��d��h�#���${�DUǼ�����w�
H�3Ꞿ�pdجJ�)�87��~��7/IG�d�RuI������<��s��;v9$k;���v�����/��y�	a�Q�@�(��ˬҋ[�[�ڳW�KjJ��m�:z!�Y�n-�k�����FX�mn`�9Z��h�%����C��Z7�kc�����D�#���ض��ٷkB�*�2�Զ�D��4�yJs�
�5�{E�
�D�"&Q>D��q;��:uI��{��,[��v�qa'�XZ2=�{<$��s�Y�Ei��x����}���c�'Op��k4@�Ԗ�4Ҍb˶��a��Gm��+����o���~��y�t�X�����r/�y��Ǐ��w'�/Q!/|_M|�9oշ�qHfJ1
D�;Z�tv���>�|C��n�6!p����������� _o}�\T�"�K����6�����[Q�.7����
�¿����>�S��t�,NWd�T�i�T�zz�`B�Y��zv����u�:���]^P���8u����}7�w{�=��[M6�0���ݳ���*�B HY���^s}\��.���q���αF"AG�	�&`�Q���nf�fK�Hˣ�T `�bܼ�1^�K{�%��@�q���T*��ڿs�����^�r��[Gu�}�>Da��K�V�?wY�V䆝'El�ǜ��-�]���}�&�r�!��F�B����}�$e$�iF}*�91�S���D�J(��g��B���2��-�{wV(�VcU󇎴���tL<i��M�W7�d]&��a#{[
L�w�9�]�q���֫$�Y�2��\�N�opq�+��З�DD�F���Ԥ���NZeKb�ԍ���ǵ�Wv�u���bB!7���koޫ�����	�r��@�eSh���p��B1����>����o5�C��������	?d�U��*�^���	�H۪*������O^z	Hx���;k�w�=�z�+9���+usӓ�P��e.���S,kn@��bcL<�֊:��R�r��T6.e��8翺g}�MJ�}*R��V���"�v�\�秮��W���o'���믪g������������V}�Kо.^�ʯ�}]y1���t�� k��7?��%12"bJ���:�M�}.���dߝOkt1�~S�&�*�^�+�6 P�lE�f�f�o]����E�ɡ{ch����؊��L`�'Q}w�wD!AF�3���ʫ�7k��u�uc9=���4/�Y/���$}�8�q~���<��ޒa��;��ͮ�<��&utV½�skUm%=�+^ӾU�|ړaܤ�{�����m�|�ۦ?ok�0�q1kj*3Tn��s����w)Ў�ßx~�#��"Y��q-�Z��	�����R��e��/��V��cX���!Hq*&��.(vQ�F.1��`����{��������ť�;�"ᇄjBOf��ܘ^*E`�譌]�n%�帥g:N�r�B�FDFM�kx�V���	)��,����އ]����_��ѓ�kFԜ���*Q�'A�u{��{���3}�����"���18�8��_PᏏ\�>�FE������z���>'{���.#�{^�4gn��i���1��V}�4��{�7�=:���dC�K������7�&�H%�y�c���T��&#�&i�.�{u@����Gki_���q]��I�����'���{G"�B�qF�_i�{j� �{A/T�:���6�+;��CE��!�}�*I�7[}y*ZB`M�r̩ۨov�L$�n�ב��雪ل"4���̵�޻���>�����͛�X��s���^�e�����o��C���gn?c;����`�ZS�6������6q���p��r�Cԡ��k�<���땡��qyKl��l�GTD`����FkX#��Xy����Y�-P䰳
��+,���S}N�e<�Uם����9�/��&�һ;U�9诮�ۋ�/sN*��>�sZ"ga����6}�{:\$���x*h�u�H7�nvP�3�75y�T��G��G"��9�] }ǳ�b�ʍ&��Ǝ�K��U�@�ūx���e��X�A�v*��Qjbo�y��H�,��݄ka	������htռ�m�3]�;q;�ʒn�a���<�'&�*�y��5 ���,(��5չ���ӮA��THUx���_N7U���j2I��1E�W9���N�T�C��|58�/}�K@�n��$���D)&z��Uk0��E7��F>UN wm͘y��(�j�/�bP�&6�&m���j����X�;77����ݼ��H�.2t���?��峇'��Q�u���ܱEZ�S���G+�<K�x����.��N�|��O:u���P!��Y�eA��e�Ɖ��B�K���eݽn��Çs��j�38���J�K+cwEn1��`\Q�U��sSn�N1�z�q��+Df����іIr�BƮcn$&�)�\�9���X�vK�P����d��	;zhU��)T�k��t�˞���3;y� �cT)������Ց�z��@P�&-RP�g��M��(�8�!s:M�	�;�R��s�pb�b��ʣt2�Ur�u�/���q
�/��Q)�@��u�����6�{���B������H@�gJR�誱N.��	���@�
ٞ#�q{�F25��O�oy��=�ӵ�̑�IM��5iw���{g� ~�����U*������c_��L�` �R�ٳ䗓# ����������=���|�� B ;�9�-��;��B�����h&�mcͫǓ�����D��O'�}��=||��b��g�Djh4�(�U|�el���V�)�e�4Zf�\�� �[��xz<	t @���734ԡ�N��L���9�s�&;�t$��!�=����N��ѵ]X�~�"b��EIJbW.VQ������7ğ]���z�_uK�-:}�S¾T�#���:����R��ST�^�95�bkilN�q_�� ���U���_g8���[SD�e6'-�;��=	1.�^|>�_զ�۝Ƌ�N��%=[q]ݚ38!B�>{��r<N|# ��{1�p�vnu�+���W�w׃joUW���>�S{F=��m�R����c�I����n�~�7 k,��ܜ3�!���kd4clL���En��βy�8ӿ���m?h�|I��NK2�q�
��T��*$t������$��\�(��It����4�8�������a@�c[��i��z�qWm���O���le�#�Z��r�N�A
1J*BL��R�2�����6�m�G_+�/�� �^�������Xv&��i�*`�Q)��7-wg�=Gҹ����뿮[9p�v�}�?��YWO��PD�������Q��>�������˿B^Z T+ "L#�:~��S��CJd���J�	�x>�{��G�:���=��������r�����q{���'#���sUUM/9�M�Ω��rrz�~Iw� ���?V����;��;!ß���W�z ��w��ʚ�SR=F���{&�h O���1	/v�#Ǘ���zy����������8��uBڜ�/�hajR�&͔F1�՘�-ly����n֮��I�/`vce�!�a@1a���n
�.4z������ٱ��-�OTn���W���\��s�ˢ��u!�fk�
�����%�ī[�\���F�!��͗h�T:�q�	�c]q\eM.�4u��������[�%�%��Ֆ�����[l��m(ih%��
 ��Be�"'��eL��_�ҋ��S��YQ��V4�:-�����������)a�l�V1/g���\�`b�a��Wy{a�{���[�sŔ�ر�ۗ�7S��ǈ/mgkƓ<�\��VjU&�?xYWP�DϦH�)��K��ͺ����nW����>�������r�T�r�����O=��$Woöp}=Y?Kz�w���-� �> �3���Ͽ7�JWR�:�Z��;Ϟ{���5��{���P.��������v�>��*��L����9��/,��y�}������:y�s}�.����B
_f���z���]F:���.Z%�+�y99u��s�G��$�|�>f�ߟo�Y��ӛ䕯//�K%��S��ק�-Ǎ���s8��v�B���U��s�cY����'JTVb�k�/��~�����K��;���c5K�_�>�>-o:�����Y�((^Q&�����;��~��fz|3�v���<�&Qǖ��Y��̟�$iw1g���
���ޜ�І�14��۩�R�+!��DsN�f��t�,�:����q�|Y���K_��ޝ^��'�1d�9�o};Q[&j�y��"U{��nu�p�����߼"<	��v��HDTB�	HJT����vX}.�wb���& o=�vv���x�9�[G�S$�橎�e��y��%l@@$	g��+��}����Ǔ�����@��7ǯf���h%�S%K�4�_y��5d�s���  �G������[1�ˍ����c9!l�s���`���d�٠��ٻ�p�j�p>�vu˪{'=|��{m>3P�.��ם~c�;�l5;S�����\���� ��폾g��U���$,@��D�����cq����  �O]s��}s��4S�|�ϼ�$��q��� %ADx�1'����x:��w46��޺2�7q{��ƕ^��M@��	A� m'j��Ɉ�C�F��4EJ�� Y�GE��7�on!�~��2�?a=xzk��x�B�9��4��d��������{�[;�x-x�����k�6�UCR���͙�6f�P��>��;<��.��[�}5��e���*c�Kt�u�?Dz���3��qYn��~�N�g0�~�0G)H![�ܯ��=��i9����3z���tW|�Axg�-��Yoi}���s6�_g���ݡI��]Kj�2��m���LiR�&�Ě�k[v�cif�a*7�d�6��]�G�H�}2��.YX����6��u��vޯ(^�D @�{;����^��g�~��%M6���n�������&R'HCz{�t��z�~W[|�{����4} pN|�������v��}��^a�Y{�˭m��,�No3�yo����Q��91���R��$���o��?�H �dlfR�x��?u�v���{n��d�d�zN�Qq_FῩ	H�$2Hd�=�>���2�!���)ܳl0Wv]Lv �f7����:�[��Ns����o^T;��;�������{`zP���y�7;}s��) }�mf\���Qg�$��O��깎��f�Ҫ����eg>����^��GsG�����W�O'�%�}�-�?! �����WC�V�gK��,�c����魻A�\�!�O�II�]�Rݻ.��]�ۧ�rW���V^>�0���.����L@!Y���!�����i� D	P��DJq�����r}	u�"9ɧ���~�vo<���,+�(�] O���-��@U!Km7MW���c�c1��{>K�@�	�����﮶�o�OO�%�v�2ۧU��?B��! ǿ�3�^��Fg�WN����>�χ#�|�����)�����c�1>B`�N�侞�����^���~�O�c�[V�Y��E���S��9�FEBJ�Eȶ����QvMS�"3�2M��wY����;��4���}ߟ��3�������=]hge
�rW$p�Fy��`hD�In�:R�scp����e��9MWZ�v��ˡ��(=GT��3���[n�������u�8�6�M�E2�S�3�[=r;�zv=��5�Mh�+m��;�ޜ�D� ���14�f������L��KI4��ip<)��ūv�5X��Iٌ�I>����`c�D�3?:��DԄ�h���a+v(J��Gb�K��-��x���ˀη��gҜ�NXS!K���L
��_<�]~���.m�I���WQ�����%�u�rBG`%Ιv������w�<_s�G}�혈%L�O_)|6����O��Z��W�����?|�g�>�'�__�˝5ɶVe�뵙]�K��	^��k�O=y=�<}���[^Ig�$�V���J�C��L���=�]���3������<�"�����>���{����Tw�	�ceK	c�e��F)�A�+�痯{�����4(�ލ�9��|���c�������#u5R�in�qum�\әͿDz� �FZ���Q������O��:]��h��e��a"�%#3<�f��`�Y��lŃ�F3+6�Ha
�T�=��w�}�u�M,�`T�uG��}NӮ����Η
� }� y;��sϳ��WI����Km�uF�N�|[u��,��Pk�����N@�-��Ǒ:l�σ}]��g�C�H �^c�Ub� 
>�>ݛz�g�B|�
VGf)QEP�H]t�0�6��Q**�mO�b��E��X�Q�l�"K�yhs#O'�� �`}X�k�n�N{-��1����O<����Ω�s��}�B"�>߳{�UӖ�m�MT�7O�{��p��'��sg[�E,B K_ټ�)��
�|�[����HN�R�2\�� �@�k*���!�o�˞�Bs��y�B�� ���z�>�p���ET�S�嶊m��m��9_qoϾ��LY��<ͷ�_�Y�Y�g�g�Q��V��r��M���΍Jؕ,�	���V��m�[gE��b9�O� ���ڷT]D���{�羬uY�_rŕ��򺼔yxI  $����z�����k��&�6S�֩ؽ���I${*�W��[��޹}]��'�'���U��E|&e# �����<���p�[��>��wy����i ��\Rc�R
>rf�p��my�K�}��B	���>�Ђ=���Xg�@%_.�i�z>r�į�;=%p<�Cz�y����˅�pnv)�����8�Y�\���a�1Q2�S��H$� �)�.�;��¶K�Q!	Q����fS�B^Q����g+��U潼gsO�w���PY�d��^��ʬ��J&aJ���mN��[c��q����b{.~�������xs�IB��]0�k�UU`��hm�l�fH�Q��/6*����r~��뾥���.U-\����u�^�6_s_+�̷���v�!��V�g����{B�T��i�m����;䗢3��=����S����;��]���N��zߥ@� ����������:�ica��S�^���^�u��v{|O%I���B��55M����S
�	Q$fWw��[�������������Ovm�z��#�C���]p����tx#�Q��S&2 |$T�D�,ͯd*#�O�����\��ށ�� 3��v��R�sQgk�Rr+�%��k^�*R�٨Q��w,����w��6ЃA���H�Z�&���~\X��?~�_ǡ�fB0rR)H@�I�O�n%��xG�$�|����\9�º��٬�G_���fz6)��}�5<Q��%F%���3�%V��f���?}����ڹ��]ۅ���]=/��ml�r*���f|�x���ӕ��3�u��k����4L�%���ʷ�/�/C! A��{�R���R����.�)�� Q�H��۠y��m�Si�4v{���?����jw���#�(�|'~���G�u���s���xS�����9����D6C�K�پ����y��S��on�_��%1�Dy�-�/�M�T
�s��Y�]�ߔ/-! ^����[o|�Y�gӵ,l�\��N����f��+,�vNhD`�� ��&rks�)�q��L���ܻR�Ƚ���ܑ>�Μ�g����h�f{��g^0��~����];�f�^�U�n�l7�j������j�EU9�
��;�9�W�&�ǿ��}�_i��jr\���&����nUG�:	|wdg���Ky�=��x%#����ڸ��y޾�L�;Nv��e��﻽Nm��
�=�|=@7����~Yjy��x��tFG���]�TGF�l����ytR�j.�fso��l`�q�NN��}Z��ԋ��뤫�9���Vs��	�sg�c��.
�2����yf�Sa�W'��[��z��j���ɮЦw�G��]P�L����ʳg�J|wN��&����� /���a�;K��ˎ����:�����\k��j�5��N�$^V�UP�#V���Ι̞�b�;��_J�t����
[q��=�ձC&AL9�9"qbNZ�s�u=���K�':=�zQ�����ȥio���ظߢr�G	��<"1Y[�) �}B���2,k�7[X��M��UP)�]F�u��y�X�N�[k�i����,D���Y��t�m[�0�.�&[�qc��{��XL�m�Js�f���n�T���Y��*�}��%e��,Nh��r��TFO%������ђ�{��]`��ʁ*�	�'x9ȋ��w:��Wg�����N���7�C.���oZ�m����m��)1h=�ًM:��.�j�B�����^=_s[�/�N�_���g�C�~���o�sgp�U���9�s0)��
�'r���W&�@��6�z�"����;o�szx-0�`���rVL���q�Y���ީ�!YS�����a$�wk;i��..���6�;���=�/k]�{=fx{�a#*�a�m�Jᘪ�F���pA=��2-�_$�][t�)+-��ڑ��^]:#���;]����P4fo�6y�&8,e8����:;s�F�o�x���S�4dјfa���:�t�<�e�pKmA٬k7k���p=���ZB��@�e܋u�ZL�:�`���Kh),t���۠�^�6��md��կ*��O���A���'Lt�o;Vm{I���Վ�fj�,mQ��	����c] �ѸT�{a3�ϡw^�[�11��M����F�ְm�l��Mc�B��/#
z�1m9p��6_\��D�v�#a�.Nպۘ�h�4��h�6�\�kV魁��
K-m��VZ�V-Jq���6av�&*ʚ�9˅2�1Q�=t��,-a6�j��ƺ��d�3p�s����Kk8ƶ�rTk)1,��5���[AҦv�R��ʭ�$�V�0�㧕ѻv�f������qY��@�4��C���R5�\��f�l�^�v���0P�n^s���+Q���؇T�9���9�8ʚ0,�1�T(V�u�8�����I��B �wmf�YǍpr���]2��.�%&3����c��m�o!ƍ�/-�sT��Ԁ-�/��c���a��o����nb6��+��լfNikG�]�u͠w@g��кu��w]x�k��5��q�ݫ��]5���tl�/I�QҪ�U,]�ۄ�J�Yw�欔<���|�i�θr�Lka���9����z:]������ܳ�8�c&c��,�.�汹���ee�CR8ԡk[tMZW����>�q�i���WP����h���n{l#�)��p�ž��G��氠��}tt.;�3�O���D]�.�,΄��ͷY5�S��l�\t�s��v��}��a�����-�Ξ�b]��k�+lV$ѕU��s�K�D�D���`�š�f�R��+2���+�VI�.�-�{�w%�k��=(�Q�ov�}�E�oi~�D�Ƭt������q�������/��(��]���ξ�m'%ާ�p�:�˴�ӹU�c7�L\�g.�����\���O��B߉��s�欶��-�?�F/{ۻ���}�=x��
��Y(Nc#f��湖�߰������ 4%*{�;o����eO³����a6z�'̕уX�{���8Y垻4l�f#[��Ő��[L�֌���w������RB��S��n5�� McB��p�.9�g-�����՝������s�Hw�;�>�oV���<�S&�=�?v�u<O��w/�ny\HuCiv����@�9*wvmڭXuFfF��]<yBe��yðH�qBX���tb����AQ{)&Ǔ�t/z4(���H�W]�Y�|}������ӹ*=����+;�{�3���E+D��wnFkU����0�S�����?+�>�B;~{���*Q��{W}<��Q^����:f��}رO���g"�:h��ڪCJΤxv��t�\1����ߝ�Q�>S�o}r�|��~�b�8�6�8j5��A�wkXA�Ǵ5��KrTT������μ{�i��6�3tE��8�
Ů�����qP�� ���t-ϗ�Dux�����H�{D��X�s���ur�t�JZ�%D�EqF�h�d���n˛�WX�j�e],�q�e�m+,Z9u�ډY���m�,�X8|�x���Vk�����A������t&�7hsőѯTivɥ�[�9t��tQj�AsZ���m1,[%4�0�%�T˪L���-heh̻Km�c0p�b�Ƃ�[u���E�Z�n���mw&�냹���ڷ(�k��fJ�Q�N1����^J�u��u�J��S�]����1������'=^�Zf����p"�Md�cj���
T}��W�����O�K�n�(��Ѷ��K�2��a���.ɮb��D�ӓ��e�:T�dH�L̜Y;/���S��ڬsl_�<� ���=������)9)�LLB�[���{GI>�pc��]y�\:]c��Z~���|H���Q$�L��2>�|���N�Ӌ�����ڮ��9^}��e�k��pu�l���9L�u��~��O�7�g_޳�v{Fӎ���<G��p����WT��q�M2h��Y=��w��z#�8B�=�|����'Lu|�6�C�������:K=~y��L�����ݮ�{��	�W�J뮉F%�4����󯿳O��n�Z���Y[���su�kj�����t A�Wo�z�o�>�u(	()B*}	L�N�]����7�\��P(M�[�&2(�9�+κ�'��(��i��A)z�����(^���{��=�x�nX��K�*��dUF�ѱ�,�}i۝��$]ب+v�Y#Z��95;�wv`�����^C��[+8i����{q�x'�w�tc�x�U�99�涢v桱�������R�4uh�S4鳷���t֭�Z�v~�O������읽��7��}.�ۗ2Rne���OBU�@%���zo
［A�33���>��"�3���^��1�
�%1���}S�}����.! {�[���^�vs���R��w�9���	�n3v�5h7Q��B:ZZ�K�l&�ĶMaXͫ��R�gÝ�S��'}�&WPW ���5﹟k����^m�x�:u�����$��M.���.�zw��J&�r�UUZ<{=ό�z#Й�۟��k>���u�؝iӚ��{�a ���;�\>����%J�#����Cʭ'j����p�<��ې{c��G��Q�T
����GH}�B��#Ï����L-�^��p�� g1�yDin�F('6�9̫�mUآ��{P���uk�K�&�Q� ���H�v���7�mm��	�p��t��|@�]�[mN������'�"JeHۜ��з�B��yz�����4����;�x�;�K��ʛ�}=�Hn��� �H�I ��r_߲�a#ǻ���}S�mk�:��z4|=Q�~V�c]kc/5WY��gX�*ݦ���W��˚kR�T�J�Q��$����#��2�ʉ�X���/���j6�5u.v*uӏ��Dv���{ܹzm��jT����74�&�F�l�<��xy�2A ����X߁�>8bw���Ep۾�6,��� %*4�{�GjfO��N��uL��l�t����4��7~���_�R� Vi�>�ik�:X�9�;�y8/��U��S)ӕ3L��=Q�F�;ɿ3Zz���#�6G7�5Ƌ? Ӿ������uε��궉���R�P��+�Ϝ@��]�i�빹jȅ�o �ܭq�g����g����m'��?6c���(�v��$�oL��td�i�z�ln�
��I��z�'�@�^#�e�����^��Z]�E|<#���<U����Y�[R�P1Զ�\���k�xZ�FyA	+���ݕ���_Ş<tӪ�]�Y�� υ��T��T���]=c76�����mu&b$�e��]Yh�M.�t�U��uUP�Q4�֜49)�o�zX����f��ŧ�ot|�)JD�x_t�o�-tL�����l��L�0��f��da
u�~��G�b��U�N�I.���iG��qޓ�����t����@���:�(>=��&�Va���V�T}�)�! ��b��'���|��\l�l���)�J���W��=B���L߾�Z�Y����"(�-�2C? @� ���o��K4�k_��VKS%L�کnmif,��;���Q2����9Zp�����.Ӆ��|4f��� 6�t}�}J��%{�e��lyj%�����l�2ԃ�>^�������)@�E����$lͮ���@q�4!�w��e�E��5�
@����  7.ܒySl���Ms��	��T���rL��6��u���{]s�L�/�o�_I�,k�#\r����̻e�&f�0[�Z+��Xp�k�Nk��v��<���KP�^������< :3E+-�.V��,��lj]�ק�>N����3A�.kH]kL;G*9pF�N�n��a�����O�����/�����\p�	�3��r�0����j>�����֞CS�	쏏c�[�S��Җ�[�l^��w([rJ3p�mE�g�Zs-���q������9~��s����3���f]*f��Z\�Z�>��>��櫯�%%�|I��D��KZ3��/�Ru!M:M���V}?��ü�*J@�	Y'�=��v�p��x��zgS8t�_FF���{�A�@�"��˷��d�T�Jt77��Nzo7�6���")�Mq��Kϼ��zE<�2ŇU���ͷ��)̴�̺�]5k
3Хi��$%$H���]��Ed���L����V���� ��ӻ�k�X��}��@K%%��4�.���}��9�J/��+�4�z?y��8+��&���ϒ^����:�l,9���l�%,���aV���A��6���w~������;ŹE�rl߽�tGN��z���8K�+f֖a�y���E��<qP���+͞
�Uf�ە%6�T�e����߇�����-x�q�(�d=�g���]��{exv-#P�S�1��Xۚ�ۿY @@�"kW��>�C-#�}9��k�l*�k^,.�g/kc�g14��T��a��uZ�f�nfݪ��̚��һ��w��3s�UU�4^��}�#�M޺��D2(���`�k���xG�����O�|K���3N�j֔ib��
0V}[�W�	�Q)t��������|��]x�ӆ	�eL�-�	br�Mޖa����������o=O%�.�u�h�G��GGg�K喾#NE�� ���H��)L��$a����-}��$E��/o|�}�4�G��d������T͐�U����� �c��4ӷmA��F��^��&\lZݮy����ޘ⛳XX. E�خi�)��69�sz+4�K鿤Pf��}�,�gԖ.xk���?Fn������//'�Z��U-ԁ4�Zӆ��Kߟ�'
-����}�~,XY��S�Y��o&֏�IT1K�i+$5����77755-�~,�/����zX��W��@�#��G�F#�|��A�H��<@l;��'�i�].2.����s�UWT2Y��gn
�ً�pC2��^�̫�]/���<�j��d33R�J�)5T=p�%~��6ս���c����!��� 	�v���'zR��^��~��3g1�H�%�:{�r*�E�����J��N�n�
yB���K���yU��?|������0p��Iy}�Nr� t�*R����o��	�jW�j��D�:����3ۼӒi��^���mO}��
_}��+#�꧜���ܾ�u��嘺�3e�0^(
]�o�Vh4�4�Ҧ�=��/�w��{�����u���Aj+^N�>p����_�;N�|����]��������Q���S�F�Գg��t�UUM��f�q��xz!h�tR�s}ϫ��k���aW++6��R��B���ё>�WĺS!,�e��X�9z�@�0��{�֔y"i�No�7�.~�U�Ň�U+�2Tΰ�jj���dQk�#�C>������*��H�uř)�.l�8�^,=T�9��`����#��N׶� ������@Yn���u)$�x(1P�#�O���C�'t���Ƚ��XĳZ���uZՖD,ݠ{/c0��.t�a�!�N��VV��\�(�˶�s��A#���޼dA�D���Q"B2�3ô�3�s�Zh��� ���O�9�mEq6�||n��w����w��8/%�w���[w&�d���\w���϶ڝ���'Bؗ#3�m���w{}��ծ�n�{}�(�o����ళ����\0�u����B��EB�᥉��U�f�t�U�S4'T:NS)��,XYY��Z�Ѕ� ���wܛ[������f�{{��H��	#�Zt|�߆MT�ۦ��_���~=�N�XQ�	;�����y'(B�|g�~�ӂ����ܫ�vxvy�gF��������xc�=�hV� @��u�V^�lb��y^z~�5o>�98?DL+ �������3O��?�UR��J]��zY����roN˯BN"$ᾯSӣ$�&�}����>�o�b�|v=����=����B.�rp)��L|߰�qD#DT�-�7�yܺ�"�����ip��r���΁�����<�=-�m�9m�MH�ټe�FƻV�\�䆤�ֶ��F�uZf5�u	��a3���VkeͅR���(Mh9�R�����*7HJ�bS��cl[�8e�-�Z�8���ˋ�������)�-�b�z�:780�8��.n�{B�c[���X�"Y�9��ƛ�g���*e�VrcGtӚ��e0JT�>yJb���|c�jR��Q��ow��׷�p������@�Pw=0·ulfi��fr'�\32�n��t��j�p���_��4���K�l.+��\�]3MdZ��b&"������' �}wkS�s"m������bÆ�7��i�GM�>���,�����B�
��E�o�ɽ����f�������NI�W��3_5�7|�p� �Y�|/_ަ�ƥ�a�����Dj����o!�����ѝ3_��D���hS7kFi��w��N�o~�ފ���H ��w��*4�������>^mT���j]T�:n�D" ^|�+��8��˘&c���k
��%0��tS��]��\E�2P_ �2bfTD�Md �ҝ��z+0VW|������
4�e���K0L��~�ӂ�ʇ�K*}K�J�le����4���BQ�J��jMcn�-Z�+u��W�������|J�;�ݛn��{�~Ϗ[�]�h��:�|雷�gs���%,<O�8D=�b�t�\���j�����JdDA��C�Ɏ�:��k>�;�v��'(�7|�2�z���d��#�A�����J�� @�$
/�Iw3'O�grӝ�Z�Y�S{8D
�*6P+�����D�_>u��C�]]2q�_�Ӹ�lc�yGTfa���E<�D�0aگ��ߢ5 #O�D�~ڼ���z�EW8oӿ=��3<�R�(Bq�=߉)MP�e:�sUMߋ4��{�xp�Θ�T�_{��{�����nli�\p]�z�њ.U��I5��)t��_!� @Y��c/�ao�3ξ��Ň��=�^�0�$B�`���~�_��HN�ʂSmʦ屹��w7�kK0��$$��o���/7��̋�ͫ�
�,�� �{��*���1m���wW�#l�f���m*��\W\5Ÿ�~I'�O8��4�e�*\�������Ϗ߻Ϊ�Gy�j��$37��د�	$�G����W=|��K<p�s��S	L����s
0��^o&��DD�����{�5~>2��j�d�.�ߪ��Lr|?�;�%��z��ګ:�ï�S�Qf��}j�/����M���=���R/�s�/�w�k�Z����%`�\W��]���N��}�wب&v���؃��������	w&s�fs�3�6�o�E������	�Q��KQ2P���3sv�s��TS}�8��}�Z��I�|���n��W��&q+.7V��ɝW�UFEht�ά��g$�1��c�8W x��-yd�s�%0���07oq��d:S7��4��؍gG4��􍬣����Ə��߻i���1F�����OÁ�A!qy���rf�h���4�Ví6g[ɻc�a�������41Ur7s����6rF�廁˩�j�m�`��H݃�XzE�;���K���ru���il���ژ��t���Wܮ6�'3f����{�3�e-��fg[��y1y8[?�)���I�g���/��e^q�E���������j|p��s�j�bp�z/�_R�*LL\�k�ݥ
i����LK��4z�����/���O��8����i�qR'>��j�Qקr��UEsGD��P%(U?y�����9�,��ϛ\P-�p���h�F�LvP�7�Qި�8�ls냛o��=?���o�z-U��Q���A�����d��ʺ7�]b�v#��1��w����u� �N��L� �_�*��>ZCѮ��l�u#�.�o�c��mM9w����˸��Jg-�����M8f�J�7������L`\�<�zgc]��Y��ѓ���Ӷ5��iK���8���O9�}�5�܉���v!l�����`�&�Q��ؽ�.qR����ۈMd^�5���b&3�9��P��S�J�>�!~�����w���l�گ\�RkL�q|e���+b�)$:L��+y���׹Tr���j1�ޜ���Uz�{�\\r�������uGN�E�ò���ANb�#!$I%����5
���vz�K��$���2����
0X��{���v�-@��^�z���z�w�+�>[�4�76,Q�E?��z/x���v����Ӳ�F�.�t����7ء�154Z�'��Ҕ�L��B��{	J�jJ2��\�de&�����>�	�5Q���Fi횷#�F����+�7�,�w���txc�%���t��Opv̯n��P
иr�E�\�{�I�7cU���$W�(ǧn�����C�13T�̅U�f�y���Tu	̐H����+��d�@�g`�T�3�Dԧ*��5���2�\U�v�UQ=��"�^�J����x�ow[��m��ד�*:�%��:��\�*���chLok����hg���$p~��#��gD�oV�Y睷�޾i) ���8ӏ����]w<�I�QE]eU�Ήn�سw���l�8Ӎ�>�j-כ;���[��
��ꔜt���>#�ZqS�d��e��xl���4,CFl�3Ӌ��b�&�nX��}�;xWUf�������×	u<P[�q�qW؂�Vt]ʝ�o�<�{��ða\�λ���{?x����JrZ��G����a���vT���z��(����u7]��bw2q��u �N�oEZ�eǉ�6R�«.q��b/���4őj��_{4����}�ʤ����1 JJ0��x�ag�:}���/�Z�`�ReL��P���Jb(@�G�MiF���b�4i��m��|l����>��d�o��P���r�P�mRi�j֔d*!>�,�֤��&>�5��4v+�qYV��a��L�,�M|=B8�Kԍf������:F]�M�N�ԭ{{uڲ�ݩ�c�q�iH�����s�E�n�pі_}�����;���������\��#� K�I<p�^ߝ�g�'��Y��Ue�u�w_�;�ò�����DD3N�z���|-Ͼ�8,�旁9�(���#����j�}B��TJ�D4q�Y�zy)<{���xQ_zT/�
�#��/����{��a񕼪�UR"��T6�2��~��P�H# O_=*������p��ņ}�rz��Ozj���sb��*��������K��(�Zr�ۚUط�xI��;J�l����k18��*o�����5݋_�ih�k���gC����e�7�c��G��D���d~A��3	��-T8�IV����A�3w���� 9Y���G��uG?����M�M7�h�=^���a}��8Q�+���Tic�zZݖi�|�W���1߳�����=vk�ct�G5e��YQ�H>����X�=�2�t������g9��F�r�X�TDJ�6F/��E����p��I��w�9}�CV��!x_}5�ӆ�y�tA��
!�w�f�N��@���d{�p�}f�|<`�}�����(�k��x�dX_�����Q+"���7}Eq�	l����M��K7'����,2c�Mf}�zY]�$�B� ^0��]���%�3�r��Re���
!SNiK���>(�@�/���=W�힓�}ɼ6�5_MGs�.1��=(��ri��<"�tU���x�����W�a��	J� J<��+G�(��%��͖Ew�k�����k��Y��} ��㱱&>D�@<�Ȼ3[�~�1Qç�]
�I��;44�z%��Rf6�ϔ��A]�2J�����7Mlq讪�]���1�K�-��
Yj�;0sY���a��.-3νɠ-#V�]�$1�BP��Eݏ����1��v����n[��Q���/$f�մ�����a�(+/vz7i�f�룭�x�κ�Ψdh��u�dcH3v����sնݷd@7_���o�;@���zF�'�v�j��QDG�'�U;W�V�m�QD��l:zܻ�p��j��z(�K���|�w{V �K���~���z���ߕ	�<��"�ca�Y��*�̖�pJUm��m/(J�Z�W"����qf���:UJ������ܽ�ZY���͹�4YS�ȯ�^����]��V|�4�Ms������T�:�Ҏ�#3~��߼�Qg�f�~�\l�p�ݖ�28a�5�]�+��T(�i�a���G�c"i�UU�B�p�sܫӂ�å^ޫ��
T�����}��Fi��;�Y��r^�5B��t�Km^����UF�����K)����if
{y�z3	�%0���H6��;�bӃ�Ѿ����D�:u-y��=������
:�BMG�=_s�4�����^9��M
�{���N����J��bTԌkS,,Zev�c�$z{p���m-�9IjR�Wkm����%��v8�*��m�:���t����RG�{+"�!���]���@��Ҥ��v��k�4�w�;�l�TR%�Q4��V`�;{�/OD{Ն^�K�W���|jւ�v��n�#Fmx�-���d����ĸ����Q�O� EB�YC�z>�и�n�s{q�<��$�{������4�g�.r���V�Б�cv�eU�7��ւ���a��$l�+��8?�3��hb_|W#���^ͭ,�|,��w���������x���*�sM�h���b�h��lފ�9��n�f��DLhD$�ܬ�w�4\?mgP����N&�SUN%�M7W��uע�I|a~}���Ō���=(�Y�r��i�a�H��'��+�i�k	�*�&M�j֌2x,ǿ;�8`���T�O�����s����جÃ�斴���6<�%Ϳ�|o?q�A�ny�rt˂�-bl�i� �T��b�����$M��T�ɥS-R�ۿ�</������,]�滽��8|^n��K @�$�m��&���Z}_z���8�
bD%��!�-��T���I�>E��~�`��j�Gb��u�tV���yϤ��O����-i��Ung^��Ҙe�b�A�enz)�?{�us���oc�����Պ<��
���2�@Om]y� T��EO��>� � ���H}���^�n�֓{r�6j�G�V�;!Mɋ-�q\V��h$�R��X��P�ai�E��5���Tz�C�����&D.���fM�D�����,�zT�0�2�d�nmn��/(W� H!|t��v�sf
�Vo��L�f�j�즊=��f8k��ĘX��^XUT�T�Km߁�a5�^,>�o�X q�/�Ug̊.~��0wVwN>���ߖR��o���k���c)�X�+�ˋ1r��M
��-�aD÷Ϝ 9{xJ&y�]K�����p�?{��\0���l�Y!b�|�w�JaG�s�=�]o=;)�ݼ�~څ�p1[�|�$���r�����%TD/�8/_���P�O��+Z����j�����ω�OLi��yZ��S�*YR�r$�ϊ��M虄u���Ӈ�P�b@D�;ɾwiQ��z���N8)gVɨt�d��	�XI��\��!o��_��;{�z.d���/U�:/B^[�~�o�����E����d@Ԍ��6��:w��j��,뭡G���o)��6��U�$Imp\*��I!	�]���3��	��o����3�f�Ļ�p�/��dS�LK/��+/:v/)�bW����+�ۙ��#�!�Pg�3���,ǵ�zY���2�J��#�S.j�_O��ߩ�3<�ah�"���B�J���꯫�"���4�Q��s�g��6 [����Wp��Iqa��Ss��&[v�8n�1bw=�ߘ�����`��ܺ��xTxV?o�ĝ,S�ݛјEf���HJ��!x��ŝ=�g&�#ŝT�V����N�5k��{��m}�o��D+K����u�ܫ^8G���x.��;[z���H�@A�g�zҩ�JuR�h)T�7�� Ǟ�X1t��ߩ賞 C ���Wʆ�?,��]W,��uUQ�Kh��n���P�p����Q�����Q�1Os�W�0:_�!m��
�����p��9��3*���;��rt�Æ�|�4��Bn��]O³x���Q;��w��Ǣkظ��ҳ_djC'fqQ�����,�"�c�Z�[7r/l)S�#Ĩ\�����$9�"HX����a����9�63����6+/R���4��յͫ���e�nrZ�-y��u�7��v��\-�V1�xRf��������.u�F�Q��كd��w=l�8ݮz�RE��I�`U��B/S�x۴�mcD������E�͓#e�rVԍ0��FVL�7i�՝k�]�H"�9�"�	�R۶K�����h	nER�|�wi
��NS�_c��{���zt&g�����/y�V���lOKZL��:�}��a's�{;<�z`K3��W����O4�69kf"T��eYm�\��:9-1V��5�v���M�����{�=����h�&�Ԓ�4ˆib���^0����
�N����?����8�t���PĦ�8B��%���i)!!ͳg���o���B��_�ok���߉��K7>�t&t�N}�^��Jb)ő�^���i�CuNo����߹7�agv�U�3ܞ��"d����i#>�s�zf 0�v���b���"��-��H��#�=��Z��d3��\kMt�����H!|^{��%�	���I���V�ן8Q���'>�<2��Z�LB=|�ѐ�}7�/K�߶�1<���_K�����*�`�cI���z��y;]��:}����v�B���{ݽ�˾wP��0$�m߂�ǅ�빼��O'����^�Ӈv����DT*D|a�������\}G��@$ap}�1z�y��O(�}���\�r������/�����R�]DH-d�� ��������4xbV�O��U��̎���Q3q�q>��d$���5��w\P�����r�C�Ph���ֆ��
��Ü�<�R�"	�pZ��f�K����} ����pϱ\Q���]�ޖ24�we�xo�G� ��$��4��M3U�S4����F�+�~�ZY��;�ۮ6v��x&���E}OEq�^��t�vS�rW�*i����G|��	��G/��~�u��7��:I��ٵ��9�
Q�{���ztf�_R�y(��	�J��&�		��^���Y��B���_�����'��&�%�8.����P�}�UI������v�n������z﮳ְ��D�Qu!�/^J����׻�����D�P�1S�������~��w�Ś:wP]}u���'�<D����xtD����ui���eS��Bxc7�O�ס7	9��'�;�b�:��~�3�cߪ�]�_RP���.0%b
(�QZ���8G�9��_%F���=¸���|(m[��tX��H-B�f�?C�?�{�wOa� ap�O�Dcp�f�eGٚ��S���i�Z���U�X>ͨDoLJFS�N���E�즳�ݳ�8���@�o����;��û�W���fֶ��a���������l��F��F��lVr��[}��0�}�f�S�T��]9��xa���Bq�G/3꾌_��z[ٌ(���n�8t�%,����{��K��'� c6T:l��ؕ�ͫ���$b��~��Q�����Tلv�noó�g=O�ݭ�.�h�q����#�7�Qg��p��it�SV<�hk+;�qX=),����&���4g=~秋��8I�zF��ȳ����{u
�3����M�\4��9�e����K����Ż����J�t��h߽��˕�C�/Å}��kOD	P���=�К�L�S#�w㆔p���}��ת�\^�S!DĚp��'�Q��z���Y���KY�&���ׁ�>��/�	>�sw�����U=�֔t�n�^����}o�>�}��#�]��}$kې � 0�!0�+� Z�Q7)���$|BA�H���PEv^���&�o�W�ȴ=�tߦi�����OI��~���[���u���7B{����S��{{�\KP�U���d 	���Xl�����'A�(��(?�A�G|���c�=	
����D�����Oљ��<+z�N{�!��UZ6l��=��.�j:�oY5Z!��A�<����d	4����!��jXۛ\,��o��^�0\6����!���}�$��%�����p�#�ɓbe	�F&+��Mj�yuxn�*�#�&W�:}�ܫ6c���^�k��*�5� ��D�����):s4ꥶ������ދ����iYO�I8�BT1{����<#/�_K\�̓f���C�����ߏ$�� !p�7�-|3
}������|.�����}	U(���ZE��6�������fu��������/���&<�ADpQ���}Wዧ�o��Y�y��\��_�~��_Ԫ� �"����D���"/W�?{V(�( �)Q��]����0D(Q@�X�W��P@O�@QV������������j���O�g�����֢�*����9����(���"�����������������G���"���?ϛ?_4g�����q��J?�0��������{�o�g���k�����q�;@�$`HFD��%!IB��!aH IXR�$dIFD��!!HIB@�!e	I��$`O�0!	R�D�� 	��%`IY��$F� HID��%dIP��$dII �!$H�$IXR��!$HXR�� @� e	YF�$ID� IXRR���%dIP�%dI`I��$`HIRD� IY�� eD�� 	 �$ I �%$I@� e		RP��$	VD�� $H��$`HD��$dHD��$RD��$%YF��%`IXD�� 	@�%$ID�� dI	BP��$	��$aIYR��D��$e		XR��% IXXB�� RXF�� IP��%%XR��  I	��!dIBD��!$H`IR���%dIHD�� $HHR��%�$ IHX �% HP��$e	XRVD��!!HdI	BD�� $HV���$%I��%�! I�� e	BD��!$HXD��!$H	D��%$IIBD��$$HI��!$HRRD�$II@�  HXRH��!�  I	BD��! H`H	@�%$HRD��!$IHR� HHdHHRP��!%	@� $IIVD�� �$!I!IFD�� %IBP��� �$ H`HHIBB��%%H%aHI�P��!� RD��%$IYBF�D��$`IR��! I��%� 	D�� YP��  HdHD��!$IH�P��%�$�"D��%�!�!�e� aHXRB��RB�BX	BXRD��% I`IH`I	R��  I!HIR��!`HIP� HdIH��%�%�$ HdIdI%`HXBP��P��!%	HP�� %	HY�D��&P���� %dHYB��%�$�$`I`I%	`HIBIX%	IB �!%`I%BD��% IP��%% H`HP��P�� � `H`H%	 HH�� H	BIYBBD�� `H%	 H	B	BD�P�D�� dHH`I% I`I IH��P��P��$ H JP���!�%�!�!� $I%RRY$HaIdIdI`H`HB�P���$� �$� �!�%�$�!� % HIBB�P����P����&�P��%�!� �% H�!�%� � %	H`H	BRP��BYB`I	BXB`H�$ H I IIBB�P��$�"�P��$�&��  He	`HYB��P��P��h@(A��B�P�@*�D@��V�V���
B�(�(A�)T��Jh�)h
��
J(((R����h* �j�h(*���d4D��QE1,�IAKKACIM4�AJSAKE@�!TД�H�KJR�4�@Ĕ�%%SAH4%3!HP44�-���)BPД�44�0�P�	HPL$@��
�Х �"�"�4#H%P4��	��б P$@����@ғ-	�+B�%+���"Ҵ� ą	BD�IBҴ�!�� PČJR-#JP*�	KCAB�#��,JR�H P	@ĉH)@R�	JDJ� P4-P,HR�B�K@����	@H�4�B4�D�H��H��R���,BD	K@Ҕ�4+JP	@д��4�IHд-
P%"P,@�H+@P4�Jб
ĢD�JD#��,BR�+H�1
D�P�	�@4-P��ʴ��(DJP4�+��)Jĭ	@�DHД�!H)H%	@�@R!J!1#��%�#H4�BP	�B�R!J�$�B��@�$�#
B�$"J@��) JȒ�$$�@Ȑ��!J��$�"JJ�$�(B��2�,�#(BH�0$@$,	 @��$��
H��$�	 H�2���@��$(@$�	 H��,	#@$�"J@�)*H�	#"H���	(H@��$!"@���$��"H�2$,	#"H$H0$��	@$,	B$�"H��,�
J$,�+"JH�$	JȒ�$)#"JȐ�)+(B��	B�2$�	)H$�)
HB�	B�2$
H��2$�(@���#JH�2$��@�2$!(@�#
BH�)	JB����"@���,�#HB�$	
JJ�$�	"J$�"B@�	 @�2���@�$	)
J��2$�@J@���H��$$	J�$�(JH��$�*p�ɉ�����*"������|o��=�����8��������?�>���TE\�y���,�_��O��_������z9�����/���~��W��#��?��/��O�UW�W��Y�^'����(���#���nn=�"����тZ�Մӟ�g����G���TEX�'���TTE_��{C�����<�'_����߁�?������QQs���~����TE_��������=�mt{������Ƹ9g�q��?�â�7ʊ��~������>�ѳǿϞo��A��W~��7���E�i8�����z�E����5��3�����~��O�?W������)����� 4��9,�������_���0߃=D  �     ���a2dɑ��4�# C �@���� h � 9�14L�2da0M4����5=$ PhM     �A�ɓ&F�L�L$����BdyFC"bd#'������5� �!���СtN���EH!�r$�(�F?��������ж�?vt$d�A��F���>.�	`"��"$`7����ϳ>�ח��Q<;�|z}~=nY�e���ʹy�����PŜ�-�аo��ڲ�´3]Њy�-N�Q���Â��IX𩃢�%���%�\h(�a*0�,q��U���U
+��wS5K��)l����Ʃ���Z̽�[ˀ�voj���]QUG�GpZ>7*����A��h#�Q���*�a��j���.X�i����6k�&���:�k[u�@։׻q���6ga��!!ܶ7���$�ES]3�d��T��IBŋN�f��X�WU�z����v
$X@�I�R�t�q�W�&����S�M���͕���0�a3�@Q�$~�V��?Nzjn�iA-J!B��-M�bdZ�a��D�q,��(fU�햘@n�6�5�q�@�i��C�3:� ҄�U�Pi���Q�gA��YaC�X����Q�  ��/�
ʽn8���J�@���/$<
�,�y�}�DV>��S
�Y6�C�ԃg�ͻ�\.��հ���Ы{���o��GG��&pvq8��)�f���S��|W��c�)V��qj���N�<�2�X�Cr�	E(6B#��(�$A�tl���ف�6lfC�:P�J-E�W�Uu�4Cү7�څa�҈��4s�8��K�
ɹP+�ո���ekL�16���rS	:�[�XA�nj��ߗ��lS+o����fq�]�q�p(}!���w9O��ߕ�PUZ������t4�oZޗY.f6�@��`|�wʛxZ�0f��ͼ]+kZolz��<A� �@��H$I| � R��`(���P�X�_�(���g������kqUb2Fp bY�B�]5U�%�M��[8e�H�PC!k"b:�8�
u\̻����p��'��w�Q!��6�E{�um1��r��Y�,X�IIc�FYq8����g�����N�V�Rj�J.M,t&A�.a��u�Ub���ކ�Y:����%�w�ک��(�0��BX����P�(:���0	�C�G�T{�s��Ð��Q3~H�ꃬ8�H@��Y��@m̀8��hm�C��!�(���c�e�������c�>���<mDdOM�����yG��ݕ��b�p�[)k5p�б|�BB� U6hĦ�X���;���������m8�b-%{���q��?���A�P�{��O�Џ@c[��HG�n{��?��޾���Oa�JXg�Yx&I�`�!�/��9'����1�Z��
�9G��sξ��5�̀�~Ӵ�j_�WҘ�y���X�u�a3���w�?c3�H��Є|�n�U!���>��P��/�I�cE	��dhy@�.�m.�j.�#�n��K���<��8j�R+!�X�X~��s�DD(H$n��.�����j1kF��A�-�HYrbz�����q��+"�g�B�p�r:��R'���h�O�=C����p���ߵ�_a�`��~%'R��P�=�̦�t�;�;M���(�F�v����m]�s��F�aD�|��8dXD�0_�/��rJ����ϙ��g.��t;�5���oGB�)}Y!`�����m���2&�>
����q��GQ����vO��/�Q��Ռlי��y���^+ڸ�f��Ň��`�C~��oSC�n!�Ͳ��n�"R�e��O��S�r��"��hK*T���d��X�' 0�ć[��2vG2��gV�ڙ�ҎP�!�2r�nk����w$S�		i�